module tapped_delay_tdc (
	output Out,
	input CLK,
    input RST,
	output [20:0] out_data,
    output reg [6:0] HEX5,
    output reg [6:0] HEX4,
    output reg [6:0] HEX3,
    output reg LED1
);

reg [1023:0] Sum2 = 4096'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
reg [1023:0] Co2 = 4096'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
reg [11:0] Sum2_hex = 0;
reg Ci = 0;
reg Selector;
reg Hit = 0;

always @(posedge CLK) begin
    if (Hit == 0) 
        Hit <= 1;
    else
        Hit <= 0;
end

reg [2:0] RSTr = 0;
always @(negedge Hit) begin
    RSTr <= {RSTr[1:0], RST};
end
wire RST_risingedge = (RSTr[2:0]==3'b001);

out_hex out_hex(.CLK(RST_risingedge), .byte_data_send(Sum2_hex[11:0]), .HEX_5(HEX5), .HEX_4(HEX4), .HEX_3(HEX3));

always @(negedge Hit) begin
    if(RST == 1) begin
        if(Sum2[1023]==0)Sum2_hex=1023;
        else if(Sum2[1022]==0)Sum2_hex=1022;
        else if(Sum2[1021]==0)Sum2_hex=1021;
        else if(Sum2[1020]==0)Sum2_hex=1020;
        else if(Sum2[1019]==0)Sum2_hex=1019;
        else if(Sum2[1018]==0)Sum2_hex=1018;
        else if(Sum2[1017]==0)Sum2_hex=1017;
        else if(Sum2[1016]==0)Sum2_hex=1016;
        else if(Sum2[1015]==0)Sum2_hex=1015;
        else if(Sum2[1014]==0)Sum2_hex=1014;
        else if(Sum2[1013]==0)Sum2_hex=1013;
        else if(Sum2[1012]==0)Sum2_hex=1012;
        else if(Sum2[1011]==0)Sum2_hex=1011;
        else if(Sum2[1010]==0)Sum2_hex=1010;
        else if(Sum2[1009]==0)Sum2_hex=1009;
        else if(Sum2[1008]==0)Sum2_hex=1008;
        else if(Sum2[1007]==0)Sum2_hex=1007;
        else if(Sum2[1006]==0)Sum2_hex=1006;
        else if(Sum2[1005]==0)Sum2_hex=1005;
        else if(Sum2[1004]==0)Sum2_hex=1004;
        else if(Sum2[1003]==0)Sum2_hex=1003;
        else if(Sum2[1002]==0)Sum2_hex=1002;
        else if(Sum2[1001]==0)Sum2_hex=1001;
        else if(Sum2[1000]==0)Sum2_hex=1000;
        else if(Sum2[999]==0)Sum2_hex=999;
        else if(Sum2[998]==0)Sum2_hex=998;
        else if(Sum2[997]==0)Sum2_hex=997;
        else if(Sum2[996]==0)Sum2_hex=996;
        else if(Sum2[995]==0)Sum2_hex=995;
        else if(Sum2[994]==0)Sum2_hex=994;
        else if(Sum2[993]==0)Sum2_hex=993;
        else if(Sum2[992]==0)Sum2_hex=992;
        else if(Sum2[991]==0)Sum2_hex=991;
        else if(Sum2[990]==0)Sum2_hex=990;
        else if(Sum2[989]==0)Sum2_hex=989;
        else if(Sum2[988]==0)Sum2_hex=988;
        else if(Sum2[987]==0)Sum2_hex=987;
        else if(Sum2[986]==0)Sum2_hex=986;
        else if(Sum2[985]==0)Sum2_hex=985;
        else if(Sum2[984]==0)Sum2_hex=984;
        else if(Sum2[983]==0)Sum2_hex=983;
        else if(Sum2[982]==0)Sum2_hex=982;
        else if(Sum2[981]==0)Sum2_hex=981;
        else if(Sum2[980]==0)Sum2_hex=980;
        else if(Sum2[979]==0)Sum2_hex=979;
        else if(Sum2[978]==0)Sum2_hex=978;
        else if(Sum2[977]==0)Sum2_hex=977;
        else if(Sum2[976]==0)Sum2_hex=976;
        else if(Sum2[975]==0)Sum2_hex=975;
        else if(Sum2[974]==0)Sum2_hex=974;
        else if(Sum2[973]==0)Sum2_hex=973;
        else if(Sum2[972]==0)Sum2_hex=972;
        else if(Sum2[971]==0)Sum2_hex=971;
        else if(Sum2[970]==0)Sum2_hex=970;
        else if(Sum2[969]==0)Sum2_hex=969;
        else if(Sum2[968]==0)Sum2_hex=968;
        else if(Sum2[967]==0)Sum2_hex=967;
        else if(Sum2[966]==0)Sum2_hex=966;
        else if(Sum2[965]==0)Sum2_hex=965;
        else if(Sum2[964]==0)Sum2_hex=964;
        else if(Sum2[963]==0)Sum2_hex=963;
        else if(Sum2[962]==0)Sum2_hex=962;
        else if(Sum2[961]==0)Sum2_hex=961;
        else if(Sum2[960]==0)Sum2_hex=960;
        else if(Sum2[959]==0)Sum2_hex=959;
        else if(Sum2[958]==0)Sum2_hex=958;
        else if(Sum2[957]==0)Sum2_hex=957;
        else if(Sum2[956]==0)Sum2_hex=956;
        else if(Sum2[955]==0)Sum2_hex=955;
        else if(Sum2[954]==0)Sum2_hex=954;
        else if(Sum2[953]==0)Sum2_hex=953;
        else if(Sum2[952]==0)Sum2_hex=952;
        else if(Sum2[951]==0)Sum2_hex=951;
        else if(Sum2[950]==0)Sum2_hex=950;
        else if(Sum2[949]==0)Sum2_hex=949;
        else if(Sum2[948]==0)Sum2_hex=948;
        else if(Sum2[947]==0)Sum2_hex=947;
        else if(Sum2[946]==0)Sum2_hex=946;
        else if(Sum2[945]==0)Sum2_hex=945;
        else if(Sum2[944]==0)Sum2_hex=944;
        else if(Sum2[943]==0)Sum2_hex=943;
        else if(Sum2[942]==0)Sum2_hex=942;
        else if(Sum2[941]==0)Sum2_hex=941;
        else if(Sum2[940]==0)Sum2_hex=940;
        else if(Sum2[939]==0)Sum2_hex=939;
        else if(Sum2[938]==0)Sum2_hex=938;
        else if(Sum2[937]==0)Sum2_hex=937;
        else if(Sum2[936]==0)Sum2_hex=936;
        else if(Sum2[935]==0)Sum2_hex=935;
        else if(Sum2[934]==0)Sum2_hex=934;
        else if(Sum2[933]==0)Sum2_hex=933;
        else if(Sum2[932]==0)Sum2_hex=932;
        else if(Sum2[931]==0)Sum2_hex=931;
        else if(Sum2[930]==0)Sum2_hex=930;
        else if(Sum2[929]==0)Sum2_hex=929;
        else if(Sum2[928]==0)Sum2_hex=928;
        else if(Sum2[927]==0)Sum2_hex=927;
        else if(Sum2[926]==0)Sum2_hex=926;
        else if(Sum2[925]==0)Sum2_hex=925;
        else if(Sum2[924]==0)Sum2_hex=924;
        else if(Sum2[923]==0)Sum2_hex=923;
        else if(Sum2[922]==0)Sum2_hex=922;
        else if(Sum2[921]==0)Sum2_hex=921;
        else if(Sum2[920]==0)Sum2_hex=920;
        else if(Sum2[919]==0)Sum2_hex=919;
        else if(Sum2[918]==0)Sum2_hex=918;
        else if(Sum2[917]==0)Sum2_hex=917;
        else if(Sum2[916]==0)Sum2_hex=916;
        else if(Sum2[915]==0)Sum2_hex=915;
        else if(Sum2[914]==0)Sum2_hex=914;
        else if(Sum2[913]==0)Sum2_hex=913;
        else if(Sum2[912]==0)Sum2_hex=912;
        else if(Sum2[911]==0)Sum2_hex=911;
        else if(Sum2[910]==0)Sum2_hex=910;
        else if(Sum2[909]==0)Sum2_hex=909;
        else if(Sum2[908]==0)Sum2_hex=908;
        else if(Sum2[907]==0)Sum2_hex=907;
        else if(Sum2[906]==0)Sum2_hex=906;
        else if(Sum2[905]==0)Sum2_hex=905;
        else if(Sum2[904]==0)Sum2_hex=904;
        else if(Sum2[903]==0)Sum2_hex=903;
        else if(Sum2[902]==0)Sum2_hex=902;
        else if(Sum2[901]==0)Sum2_hex=901;
        else if(Sum2[900]==0)Sum2_hex=900;
        else if(Sum2[899]==0)Sum2_hex=899;
        else if(Sum2[898]==0)Sum2_hex=898;
        else if(Sum2[897]==0)Sum2_hex=897;
        else if(Sum2[896]==0)Sum2_hex=896;
        else if(Sum2[895]==0)Sum2_hex=895;
        else if(Sum2[894]==0)Sum2_hex=894;
        else if(Sum2[893]==0)Sum2_hex=893;
        else if(Sum2[892]==0)Sum2_hex=892;
        else if(Sum2[891]==0)Sum2_hex=891;
        else if(Sum2[890]==0)Sum2_hex=890;
        else if(Sum2[889]==0)Sum2_hex=889;
        else if(Sum2[888]==0)Sum2_hex=888;
        else if(Sum2[887]==0)Sum2_hex=887;
        else if(Sum2[886]==0)Sum2_hex=886;
        else if(Sum2[885]==0)Sum2_hex=885;
        else if(Sum2[884]==0)Sum2_hex=884;
        else if(Sum2[883]==0)Sum2_hex=883;
        else if(Sum2[882]==0)Sum2_hex=882;
        else if(Sum2[881]==0)Sum2_hex=881;
        else if(Sum2[880]==0)Sum2_hex=880;
        else if(Sum2[879]==0)Sum2_hex=879;
        else if(Sum2[878]==0)Sum2_hex=878;
        else if(Sum2[877]==0)Sum2_hex=877;
        else if(Sum2[876]==0)Sum2_hex=876;
        else if(Sum2[875]==0)Sum2_hex=875;
        else if(Sum2[874]==0)Sum2_hex=874;
        else if(Sum2[873]==0)Sum2_hex=873;
        else if(Sum2[872]==0)Sum2_hex=872;
        else if(Sum2[871]==0)Sum2_hex=871;
        else if(Sum2[870]==0)Sum2_hex=870;
        else if(Sum2[869]==0)Sum2_hex=869;
        else if(Sum2[868]==0)Sum2_hex=868;
        else if(Sum2[867]==0)Sum2_hex=867;
        else if(Sum2[866]==0)Sum2_hex=866;
        else if(Sum2[865]==0)Sum2_hex=865;
        else if(Sum2[864]==0)Sum2_hex=864;
        else if(Sum2[863]==0)Sum2_hex=863;
        else if(Sum2[862]==0)Sum2_hex=862;
        else if(Sum2[861]==0)Sum2_hex=861;
        else if(Sum2[860]==0)Sum2_hex=860;
        else if(Sum2[859]==0)Sum2_hex=859;
        else if(Sum2[858]==0)Sum2_hex=858;
        else if(Sum2[857]==0)Sum2_hex=857;
        else if(Sum2[856]==0)Sum2_hex=856;
        else if(Sum2[855]==0)Sum2_hex=855;
        else if(Sum2[854]==0)Sum2_hex=854;
        else if(Sum2[853]==0)Sum2_hex=853;
        else if(Sum2[852]==0)Sum2_hex=852;
        else if(Sum2[851]==0)Sum2_hex=851;
        else if(Sum2[850]==0)Sum2_hex=850;
        else if(Sum2[849]==0)Sum2_hex=849;
        else if(Sum2[848]==0)Sum2_hex=848;
        else if(Sum2[847]==0)Sum2_hex=847;
        else if(Sum2[846]==0)Sum2_hex=846;
        else if(Sum2[845]==0)Sum2_hex=845;
        else if(Sum2[844]==0)Sum2_hex=844;
        else if(Sum2[843]==0)Sum2_hex=843;
        else if(Sum2[842]==0)Sum2_hex=842;
        else if(Sum2[841]==0)Sum2_hex=841;
        else if(Sum2[840]==0)Sum2_hex=840;
        else if(Sum2[839]==0)Sum2_hex=839;
        else if(Sum2[838]==0)Sum2_hex=838;
        else if(Sum2[837]==0)Sum2_hex=837;
        else if(Sum2[836]==0)Sum2_hex=836;
        else if(Sum2[835]==0)Sum2_hex=835;
        else if(Sum2[834]==0)Sum2_hex=834;
        else if(Sum2[833]==0)Sum2_hex=833;
        else if(Sum2[832]==0)Sum2_hex=832;
        else if(Sum2[831]==0)Sum2_hex=831;
        else if(Sum2[830]==0)Sum2_hex=830;
        else if(Sum2[829]==0)Sum2_hex=829;
        else if(Sum2[828]==0)Sum2_hex=828;
        else if(Sum2[827]==0)Sum2_hex=827;
        else if(Sum2[826]==0)Sum2_hex=826;
        else if(Sum2[825]==0)Sum2_hex=825;
        else if(Sum2[824]==0)Sum2_hex=824;
        else if(Sum2[823]==0)Sum2_hex=823;
        else if(Sum2[822]==0)Sum2_hex=822;
        else if(Sum2[821]==0)Sum2_hex=821;
        else if(Sum2[820]==0)Sum2_hex=820;
        else if(Sum2[819]==0)Sum2_hex=819;
        else if(Sum2[818]==0)Sum2_hex=818;
        else if(Sum2[817]==0)Sum2_hex=817;
        else if(Sum2[816]==0)Sum2_hex=816;
        else if(Sum2[815]==0)Sum2_hex=815;
        else if(Sum2[814]==0)Sum2_hex=814;
        else if(Sum2[813]==0)Sum2_hex=813;
        else if(Sum2[812]==0)Sum2_hex=812;
        else if(Sum2[811]==0)Sum2_hex=811;
        else if(Sum2[810]==0)Sum2_hex=810;
        else if(Sum2[809]==0)Sum2_hex=809;
        else if(Sum2[808]==0)Sum2_hex=808;
        else if(Sum2[807]==0)Sum2_hex=807;
        else if(Sum2[806]==0)Sum2_hex=806;
        else if(Sum2[805]==0)Sum2_hex=805;
        else if(Sum2[804]==0)Sum2_hex=804;
        else if(Sum2[803]==0)Sum2_hex=803;
        else if(Sum2[802]==0)Sum2_hex=802;
        else if(Sum2[801]==0)Sum2_hex=801;
        else if(Sum2[800]==0)Sum2_hex=800;
        else if(Sum2[799]==0)Sum2_hex=799;
        else if(Sum2[798]==0)Sum2_hex=798;
        else if(Sum2[797]==0)Sum2_hex=797;
        else if(Sum2[796]==0)Sum2_hex=796;
        else if(Sum2[795]==0)Sum2_hex=795;
        else if(Sum2[794]==0)Sum2_hex=794;
        else if(Sum2[793]==0)Sum2_hex=793;
        else if(Sum2[792]==0)Sum2_hex=792;
        else if(Sum2[791]==0)Sum2_hex=791;
        else if(Sum2[790]==0)Sum2_hex=790;
        else if(Sum2[789]==0)Sum2_hex=789;
        else if(Sum2[788]==0)Sum2_hex=788;
        else if(Sum2[787]==0)Sum2_hex=787;
        else if(Sum2[786]==0)Sum2_hex=786;
        else if(Sum2[785]==0)Sum2_hex=785;
        else if(Sum2[784]==0)Sum2_hex=784;
        else if(Sum2[783]==0)Sum2_hex=783;
        else if(Sum2[782]==0)Sum2_hex=782;
        else if(Sum2[781]==0)Sum2_hex=781;
        else if(Sum2[780]==0)Sum2_hex=780;
        else if(Sum2[779]==0)Sum2_hex=779;
        else if(Sum2[778]==0)Sum2_hex=778;
        else if(Sum2[777]==0)Sum2_hex=777;
        else if(Sum2[776]==0)Sum2_hex=776;
        else if(Sum2[775]==0)Sum2_hex=775;
        else if(Sum2[774]==0)Sum2_hex=774;
        else if(Sum2[773]==0)Sum2_hex=773;
        else if(Sum2[772]==0)Sum2_hex=772;
        else if(Sum2[771]==0)Sum2_hex=771;
        else if(Sum2[770]==0)Sum2_hex=770;
        else if(Sum2[769]==0)Sum2_hex=769;
        else if(Sum2[768]==0)Sum2_hex=768;
        else if(Sum2[767]==0)Sum2_hex=767;
        else if(Sum2[766]==0)Sum2_hex=766;
        else if(Sum2[765]==0)Sum2_hex=765;
        else if(Sum2[764]==0)Sum2_hex=764;
        else if(Sum2[763]==0)Sum2_hex=763;
        else if(Sum2[762]==0)Sum2_hex=762;
        else if(Sum2[761]==0)Sum2_hex=761;
        else if(Sum2[760]==0)Sum2_hex=760;
        else if(Sum2[759]==0)Sum2_hex=759;
        else if(Sum2[758]==0)Sum2_hex=758;
        else if(Sum2[757]==0)Sum2_hex=757;
        else if(Sum2[756]==0)Sum2_hex=756;
        else if(Sum2[755]==0)Sum2_hex=755;
        else if(Sum2[754]==0)Sum2_hex=754;
        else if(Sum2[753]==0)Sum2_hex=753;
        else if(Sum2[752]==0)Sum2_hex=752;
        else if(Sum2[751]==0)Sum2_hex=751;
        else if(Sum2[750]==0)Sum2_hex=750;
        else if(Sum2[749]==0)Sum2_hex=749;
        else if(Sum2[748]==0)Sum2_hex=748;
        else if(Sum2[747]==0)Sum2_hex=747;
        else if(Sum2[746]==0)Sum2_hex=746;
        else if(Sum2[745]==0)Sum2_hex=745;
        else if(Sum2[744]==0)Sum2_hex=744;
        else if(Sum2[743]==0)Sum2_hex=743;
        else if(Sum2[742]==0)Sum2_hex=742;
        else if(Sum2[741]==0)Sum2_hex=741;
        else if(Sum2[740]==0)Sum2_hex=740;
        else if(Sum2[739]==0)Sum2_hex=739;
        else if(Sum2[738]==0)Sum2_hex=738;
        else if(Sum2[737]==0)Sum2_hex=737;
        else if(Sum2[736]==0)Sum2_hex=736;
        else if(Sum2[735]==0)Sum2_hex=735;
        else if(Sum2[734]==0)Sum2_hex=734;
        else if(Sum2[733]==0)Sum2_hex=733;
        else if(Sum2[732]==0)Sum2_hex=732;
        else if(Sum2[731]==0)Sum2_hex=731;
        else if(Sum2[730]==0)Sum2_hex=730;
        else if(Sum2[729]==0)Sum2_hex=729;
        else if(Sum2[728]==0)Sum2_hex=728;
        else if(Sum2[727]==0)Sum2_hex=727;
        else if(Sum2[726]==0)Sum2_hex=726;
        else if(Sum2[725]==0)Sum2_hex=725;
        else if(Sum2[724]==0)Sum2_hex=724;
        else if(Sum2[723]==0)Sum2_hex=723;
        else if(Sum2[722]==0)Sum2_hex=722;
        else if(Sum2[721]==0)Sum2_hex=721;
        else if(Sum2[720]==0)Sum2_hex=720;
        else if(Sum2[719]==0)Sum2_hex=719;
        else if(Sum2[718]==0)Sum2_hex=718;
        else if(Sum2[717]==0)Sum2_hex=717;
        else if(Sum2[716]==0)Sum2_hex=716;
        else if(Sum2[715]==0)Sum2_hex=715;
        else if(Sum2[714]==0)Sum2_hex=714;
        else if(Sum2[713]==0)Sum2_hex=713;
        else if(Sum2[712]==0)Sum2_hex=712;
        else if(Sum2[711]==0)Sum2_hex=711;
        else if(Sum2[710]==0)Sum2_hex=710;
        else if(Sum2[709]==0)Sum2_hex=709;
        else if(Sum2[708]==0)Sum2_hex=708;
        else if(Sum2[707]==0)Sum2_hex=707;
        else if(Sum2[706]==0)Sum2_hex=706;
        else if(Sum2[705]==0)Sum2_hex=705;
        else if(Sum2[704]==0)Sum2_hex=704;
        else if(Sum2[703]==0)Sum2_hex=703;
        else if(Sum2[702]==0)Sum2_hex=702;
        else if(Sum2[701]==0)Sum2_hex=701;
        else if(Sum2[700]==0)Sum2_hex=700;
        else if(Sum2[699]==0)Sum2_hex=699;
        else if(Sum2[698]==0)Sum2_hex=698;
        else if(Sum2[697]==0)Sum2_hex=697;
        else if(Sum2[696]==0)Sum2_hex=696;
        else if(Sum2[695]==0)Sum2_hex=695;
        else if(Sum2[694]==0)Sum2_hex=694;
        else if(Sum2[693]==0)Sum2_hex=693;
        else if(Sum2[692]==0)Sum2_hex=692;
        else if(Sum2[691]==0)Sum2_hex=691;
        else if(Sum2[690]==0)Sum2_hex=690;
        else if(Sum2[689]==0)Sum2_hex=689;
        else if(Sum2[688]==0)Sum2_hex=688;
        else if(Sum2[687]==0)Sum2_hex=687;
        else if(Sum2[686]==0)Sum2_hex=686;
        else if(Sum2[685]==0)Sum2_hex=685;
        else if(Sum2[684]==0)Sum2_hex=684;
        else if(Sum2[683]==0)Sum2_hex=683;
        else if(Sum2[682]==0)Sum2_hex=682;
        else if(Sum2[681]==0)Sum2_hex=681;
        else if(Sum2[680]==0)Sum2_hex=680;
        else if(Sum2[679]==0)Sum2_hex=679;
        else if(Sum2[678]==0)Sum2_hex=678;
        else if(Sum2[677]==0)Sum2_hex=677;
        else if(Sum2[676]==0)Sum2_hex=676;
        else if(Sum2[675]==0)Sum2_hex=675;
        else if(Sum2[674]==0)Sum2_hex=674;
        else if(Sum2[673]==0)Sum2_hex=673;
        else if(Sum2[672]==0)Sum2_hex=672;
        else if(Sum2[671]==0)Sum2_hex=671;
        else if(Sum2[670]==0)Sum2_hex=670;
        else if(Sum2[669]==0)Sum2_hex=669;
        else if(Sum2[668]==0)Sum2_hex=668;
        else if(Sum2[667]==0)Sum2_hex=667;
        else if(Sum2[666]==0)Sum2_hex=666;
        else if(Sum2[665]==0)Sum2_hex=665;
        else if(Sum2[664]==0)Sum2_hex=664;
        else if(Sum2[663]==0)Sum2_hex=663;
        else if(Sum2[662]==0)Sum2_hex=662;
        else if(Sum2[661]==0)Sum2_hex=661;
        else if(Sum2[660]==0)Sum2_hex=660;
        else if(Sum2[659]==0)Sum2_hex=659;
        else if(Sum2[658]==0)Sum2_hex=658;
        else if(Sum2[657]==0)Sum2_hex=657;
        else if(Sum2[656]==0)Sum2_hex=656;
        else if(Sum2[655]==0)Sum2_hex=655;
        else if(Sum2[654]==0)Sum2_hex=654;
        else if(Sum2[653]==0)Sum2_hex=653;
        else if(Sum2[652]==0)Sum2_hex=652;
        else if(Sum2[651]==0)Sum2_hex=651;
        else if(Sum2[650]==0)Sum2_hex=650;
        else if(Sum2[649]==0)Sum2_hex=649;
        else if(Sum2[648]==0)Sum2_hex=648;
        else if(Sum2[647]==0)Sum2_hex=647;
        else if(Sum2[646]==0)Sum2_hex=646;
        else if(Sum2[645]==0)Sum2_hex=645;
        else if(Sum2[644]==0)Sum2_hex=644;
        else if(Sum2[643]==0)Sum2_hex=643;
        else if(Sum2[642]==0)Sum2_hex=642;
        else if(Sum2[641]==0)Sum2_hex=641;
        else if(Sum2[640]==0)Sum2_hex=640;
        else if(Sum2[639]==0)Sum2_hex=639;
        else if(Sum2[638]==0)Sum2_hex=638;
        else if(Sum2[637]==0)Sum2_hex=637;
        else if(Sum2[636]==0)Sum2_hex=636;
        else if(Sum2[635]==0)Sum2_hex=635;
        else if(Sum2[634]==0)Sum2_hex=634;
        else if(Sum2[633]==0)Sum2_hex=633;
        else if(Sum2[632]==0)Sum2_hex=632;
        else if(Sum2[631]==0)Sum2_hex=631;
        else if(Sum2[630]==0)Sum2_hex=630;
        else if(Sum2[629]==0)Sum2_hex=629;
        else if(Sum2[628]==0)Sum2_hex=628;
        else if(Sum2[627]==0)Sum2_hex=627;
        else if(Sum2[626]==0)Sum2_hex=626;
        else if(Sum2[625]==0)Sum2_hex=625;
        else if(Sum2[624]==0)Sum2_hex=624;
        else if(Sum2[623]==0)Sum2_hex=623;
        else if(Sum2[622]==0)Sum2_hex=622;
        else if(Sum2[621]==0)Sum2_hex=621;
        else if(Sum2[620]==0)Sum2_hex=620;
        else if(Sum2[619]==0)Sum2_hex=619;
        else if(Sum2[618]==0)Sum2_hex=618;
        else if(Sum2[617]==0)Sum2_hex=617;
        else if(Sum2[616]==0)Sum2_hex=616;
        else if(Sum2[615]==0)Sum2_hex=615;
        else if(Sum2[614]==0)Sum2_hex=614;
        else if(Sum2[613]==0)Sum2_hex=613;
        else if(Sum2[612]==0)Sum2_hex=612;
        else if(Sum2[611]==0)Sum2_hex=611;
        else if(Sum2[610]==0)Sum2_hex=610;
        else if(Sum2[609]==0)Sum2_hex=609;
        else if(Sum2[608]==0)Sum2_hex=608;
        else if(Sum2[607]==0)Sum2_hex=607;
        else if(Sum2[606]==0)Sum2_hex=606;
        else if(Sum2[605]==0)Sum2_hex=605;
        else if(Sum2[604]==0)Sum2_hex=604;
        else if(Sum2[603]==0)Sum2_hex=603;
        else if(Sum2[602]==0)Sum2_hex=602;
        else if(Sum2[601]==0)Sum2_hex=601;
        else if(Sum2[600]==0)Sum2_hex=600;
        else if(Sum2[599]==0)Sum2_hex=599;
        else if(Sum2[598]==0)Sum2_hex=598;
        else if(Sum2[597]==0)Sum2_hex=597;
        else if(Sum2[596]==0)Sum2_hex=596;
        else if(Sum2[595]==0)Sum2_hex=595;
        else if(Sum2[594]==0)Sum2_hex=594;
        else if(Sum2[593]==0)Sum2_hex=593;
        else if(Sum2[592]==0)Sum2_hex=592;
        else if(Sum2[591]==0)Sum2_hex=591;
        else if(Sum2[590]==0)Sum2_hex=590;
        else if(Sum2[589]==0)Sum2_hex=589;
        else if(Sum2[588]==0)Sum2_hex=588;
        else if(Sum2[587]==0)Sum2_hex=587;
        else if(Sum2[586]==0)Sum2_hex=586;
        else if(Sum2[585]==0)Sum2_hex=585;
        else if(Sum2[584]==0)Sum2_hex=584;
        else if(Sum2[583]==0)Sum2_hex=583;
        else if(Sum2[582]==0)Sum2_hex=582;
        else if(Sum2[581]==0)Sum2_hex=581;
        else if(Sum2[580]==0)Sum2_hex=580;
        else if(Sum2[579]==0)Sum2_hex=579;
        else if(Sum2[578]==0)Sum2_hex=578;
        else if(Sum2[577]==0)Sum2_hex=577;
        else if(Sum2[576]==0)Sum2_hex=576;
        else if(Sum2[575]==0)Sum2_hex=575;
        else if(Sum2[574]==0)Sum2_hex=574;
        else if(Sum2[573]==0)Sum2_hex=573;
        else if(Sum2[572]==0)Sum2_hex=572;
        else if(Sum2[571]==0)Sum2_hex=571;
        else if(Sum2[570]==0)Sum2_hex=570;
        else if(Sum2[569]==0)Sum2_hex=569;
        else if(Sum2[568]==0)Sum2_hex=568;
        else if(Sum2[567]==0)Sum2_hex=567;
        else if(Sum2[566]==0)Sum2_hex=566;
        else if(Sum2[565]==0)Sum2_hex=565;
        else if(Sum2[564]==0)Sum2_hex=564;
        else if(Sum2[563]==0)Sum2_hex=563;
        else if(Sum2[562]==0)Sum2_hex=562;
        else if(Sum2[561]==0)Sum2_hex=561;
        else if(Sum2[560]==0)Sum2_hex=560;
        else if(Sum2[559]==0)Sum2_hex=559;
        else if(Sum2[558]==0)Sum2_hex=558;
        else if(Sum2[557]==0)Sum2_hex=557;
        else if(Sum2[556]==0)Sum2_hex=556;
        else if(Sum2[555]==0)Sum2_hex=555;
        else if(Sum2[554]==0)Sum2_hex=554;
        else if(Sum2[553]==0)Sum2_hex=553;
        else if(Sum2[552]==0)Sum2_hex=552;
        else if(Sum2[551]==0)Sum2_hex=551;
        else if(Sum2[550]==0)Sum2_hex=550;
        else if(Sum2[549]==0)Sum2_hex=549;
        else if(Sum2[548]==0)Sum2_hex=548;
        else if(Sum2[547]==0)Sum2_hex=547;
        else if(Sum2[546]==0)Sum2_hex=546;
        else if(Sum2[545]==0)Sum2_hex=545;
        else if(Sum2[544]==0)Sum2_hex=544;
        else if(Sum2[543]==0)Sum2_hex=543;
        else if(Sum2[542]==0)Sum2_hex=542;
        else if(Sum2[541]==0)Sum2_hex=541;
        else if(Sum2[540]==0)Sum2_hex=540;
        else if(Sum2[539]==0)Sum2_hex=539;
        else if(Sum2[538]==0)Sum2_hex=538;
        else if(Sum2[537]==0)Sum2_hex=537;
        else if(Sum2[536]==0)Sum2_hex=536;
        else if(Sum2[535]==0)Sum2_hex=535;
        else if(Sum2[534]==0)Sum2_hex=534;
        else if(Sum2[533]==0)Sum2_hex=533;
        else if(Sum2[532]==0)Sum2_hex=532;
        else if(Sum2[531]==0)Sum2_hex=531;
        else if(Sum2[530]==0)Sum2_hex=530;
        else if(Sum2[529]==0)Sum2_hex=529;
        else if(Sum2[528]==0)Sum2_hex=528;
        else if(Sum2[527]==0)Sum2_hex=527;
        else if(Sum2[526]==0)Sum2_hex=526;
        else if(Sum2[525]==0)Sum2_hex=525;
        else if(Sum2[524]==0)Sum2_hex=524;
        else if(Sum2[523]==0)Sum2_hex=523;
        else if(Sum2[522]==0)Sum2_hex=522;
        else if(Sum2[521]==0)Sum2_hex=521;
        else if(Sum2[520]==0)Sum2_hex=520;
        else if(Sum2[519]==0)Sum2_hex=519;
        else if(Sum2[518]==0)Sum2_hex=518;
        else if(Sum2[517]==0)Sum2_hex=517;
        else if(Sum2[516]==0)Sum2_hex=516;
        else if(Sum2[515]==0)Sum2_hex=515;
        else if(Sum2[514]==0)Sum2_hex=514;
        else if(Sum2[513]==0)Sum2_hex=513;
        else if(Sum2[512]==0)Sum2_hex=512;
        else if(Sum2[511]==0)Sum2_hex=511;
        else if(Sum2[510]==0)Sum2_hex=510;
        else if(Sum2[509]==0)Sum2_hex=509;
        else if(Sum2[508]==0)Sum2_hex=508;
        else if(Sum2[507]==0)Sum2_hex=507;
        else if(Sum2[506]==0)Sum2_hex=506;
        else if(Sum2[505]==0)Sum2_hex=505;
        else if(Sum2[504]==0)Sum2_hex=504;
        else if(Sum2[503]==0)Sum2_hex=503;
        else if(Sum2[502]==0)Sum2_hex=502;
        else if(Sum2[501]==0)Sum2_hex=501;
        else if(Sum2[500]==0)Sum2_hex=500;
        else if(Sum2[499]==0)Sum2_hex=499;
        else if(Sum2[498]==0)Sum2_hex=498;
        else if(Sum2[497]==0)Sum2_hex=497;
        else if(Sum2[496]==0)Sum2_hex=496;
        else if(Sum2[495]==0)Sum2_hex=495;
        else if(Sum2[494]==0)Sum2_hex=494;
        else if(Sum2[493]==0)Sum2_hex=493;
        else if(Sum2[492]==0)Sum2_hex=492;
        else if(Sum2[491]==0)Sum2_hex=491;
        else if(Sum2[490]==0)Sum2_hex=490;
        else if(Sum2[489]==0)Sum2_hex=489;
        else if(Sum2[488]==0)Sum2_hex=488;
        else if(Sum2[487]==0)Sum2_hex=487;
        else if(Sum2[486]==0)Sum2_hex=486;
        else if(Sum2[485]==0)Sum2_hex=485;
        else if(Sum2[484]==0)Sum2_hex=484;
        else if(Sum2[483]==0)Sum2_hex=483;
        else if(Sum2[482]==0)Sum2_hex=482;
        else if(Sum2[481]==0)Sum2_hex=481;
        else if(Sum2[480]==0)Sum2_hex=480;
        else if(Sum2[479]==0)Sum2_hex=479;
        else if(Sum2[478]==0)Sum2_hex=478;
        else if(Sum2[477]==0)Sum2_hex=477;
        else if(Sum2[476]==0)Sum2_hex=476;
        else if(Sum2[475]==0)Sum2_hex=475;
        else if(Sum2[474]==0)Sum2_hex=474;
        else if(Sum2[473]==0)Sum2_hex=473;
        else if(Sum2[472]==0)Sum2_hex=472;
        else if(Sum2[471]==0)Sum2_hex=471;
        else if(Sum2[470]==0)Sum2_hex=470;
        else if(Sum2[469]==0)Sum2_hex=469;
        else if(Sum2[468]==0)Sum2_hex=468;
        else if(Sum2[467]==0)Sum2_hex=467;
        else if(Sum2[466]==0)Sum2_hex=466;
        else if(Sum2[465]==0)Sum2_hex=465;
        else if(Sum2[464]==0)Sum2_hex=464;
        else if(Sum2[463]==0)Sum2_hex=463;
        else if(Sum2[462]==0)Sum2_hex=462;
        else if(Sum2[461]==0)Sum2_hex=461;
        else if(Sum2[460]==0)Sum2_hex=460;
        else if(Sum2[459]==0)Sum2_hex=459;
        else if(Sum2[458]==0)Sum2_hex=458;
        else if(Sum2[457]==0)Sum2_hex=457;
        else if(Sum2[456]==0)Sum2_hex=456;
        else if(Sum2[455]==0)Sum2_hex=455;
        else if(Sum2[454]==0)Sum2_hex=454;
        else if(Sum2[453]==0)Sum2_hex=453;
        else if(Sum2[452]==0)Sum2_hex=452;
        else if(Sum2[451]==0)Sum2_hex=451;
        else if(Sum2[450]==0)Sum2_hex=450;
        else if(Sum2[449]==0)Sum2_hex=449;
        else if(Sum2[448]==0)Sum2_hex=448;
        else if(Sum2[447]==0)Sum2_hex=447;
        else if(Sum2[446]==0)Sum2_hex=446;
        else if(Sum2[445]==0)Sum2_hex=445;
        else if(Sum2[444]==0)Sum2_hex=444;
        else if(Sum2[443]==0)Sum2_hex=443;
        else if(Sum2[442]==0)Sum2_hex=442;
        else if(Sum2[441]==0)Sum2_hex=441;
        else if(Sum2[440]==0)Sum2_hex=440;
        else if(Sum2[439]==0)Sum2_hex=439;
        else if(Sum2[438]==0)Sum2_hex=438;
        else if(Sum2[437]==0)Sum2_hex=437;
        else if(Sum2[436]==0)Sum2_hex=436;
        else if(Sum2[435]==0)Sum2_hex=435;
        else if(Sum2[434]==0)Sum2_hex=434;
        else if(Sum2[433]==0)Sum2_hex=433;
        else if(Sum2[432]==0)Sum2_hex=432;
        else if(Sum2[431]==0)Sum2_hex=431;
        else if(Sum2[430]==0)Sum2_hex=430;
        else if(Sum2[429]==0)Sum2_hex=429;
        else if(Sum2[428]==0)Sum2_hex=428;
        else if(Sum2[427]==0)Sum2_hex=427;
        else if(Sum2[426]==0)Sum2_hex=426;
        else if(Sum2[425]==0)Sum2_hex=425;
        else if(Sum2[424]==0)Sum2_hex=424;
        else if(Sum2[423]==0)Sum2_hex=423;
        else if(Sum2[422]==0)Sum2_hex=422;
        else if(Sum2[421]==0)Sum2_hex=421;
        else if(Sum2[420]==0)Sum2_hex=420;
        else if(Sum2[419]==0)Sum2_hex=419;
        else if(Sum2[418]==0)Sum2_hex=418;
        else if(Sum2[417]==0)Sum2_hex=417;
        else if(Sum2[416]==0)Sum2_hex=416;
        else if(Sum2[415]==0)Sum2_hex=415;
        else if(Sum2[414]==0)Sum2_hex=414;
        else if(Sum2[413]==0)Sum2_hex=413;
        else if(Sum2[412]==0)Sum2_hex=412;
        else if(Sum2[411]==0)Sum2_hex=411;
        else if(Sum2[410]==0)Sum2_hex=410;
        else if(Sum2[409]==0)Sum2_hex=409;
        else if(Sum2[408]==0)Sum2_hex=408;
        else if(Sum2[407]==0)Sum2_hex=407;
        else if(Sum2[406]==0)Sum2_hex=406;
        else if(Sum2[405]==0)Sum2_hex=405;
        else if(Sum2[404]==0)Sum2_hex=404;
        else if(Sum2[403]==0)Sum2_hex=403;
        else if(Sum2[402]==0)Sum2_hex=402;
        else if(Sum2[401]==0)Sum2_hex=401;
        else if(Sum2[400]==0)Sum2_hex=400;
        else if(Sum2[399]==0)Sum2_hex=399;
        else if(Sum2[398]==0)Sum2_hex=398;
        else if(Sum2[397]==0)Sum2_hex=397;
        else if(Sum2[396]==0)Sum2_hex=396;
        else if(Sum2[395]==0)Sum2_hex=395;
        else if(Sum2[394]==0)Sum2_hex=394;
        else if(Sum2[393]==0)Sum2_hex=393;
        else if(Sum2[392]==0)Sum2_hex=392;
        else if(Sum2[391]==0)Sum2_hex=391;
        else if(Sum2[390]==0)Sum2_hex=390;
        else if(Sum2[389]==0)Sum2_hex=389;
        else if(Sum2[388]==0)Sum2_hex=388;
        else if(Sum2[387]==0)Sum2_hex=387;
        else if(Sum2[386]==0)Sum2_hex=386;
        else if(Sum2[385]==0)Sum2_hex=385;
        else if(Sum2[384]==0)Sum2_hex=384;
        else if(Sum2[383]==0)Sum2_hex=383;
        else if(Sum2[382]==0)Sum2_hex=382;
        else if(Sum2[381]==0)Sum2_hex=381;
        else if(Sum2[380]==0)Sum2_hex=380;
        else if(Sum2[379]==0)Sum2_hex=379;
        else if(Sum2[378]==0)Sum2_hex=378;
        else if(Sum2[377]==0)Sum2_hex=377;
        else if(Sum2[376]==0)Sum2_hex=376;
        else if(Sum2[375]==0)Sum2_hex=375;
        else if(Sum2[374]==0)Sum2_hex=374;
        else if(Sum2[373]==0)Sum2_hex=373;
        else if(Sum2[372]==0)Sum2_hex=372;
        else if(Sum2[371]==0)Sum2_hex=371;
        else if(Sum2[370]==0)Sum2_hex=370;
        else if(Sum2[369]==0)Sum2_hex=369;
        else if(Sum2[368]==0)Sum2_hex=368;
        else if(Sum2[367]==0)Sum2_hex=367;
        else if(Sum2[366]==0)Sum2_hex=366;
        else if(Sum2[365]==0)Sum2_hex=365;
        else if(Sum2[364]==0)Sum2_hex=364;
        else if(Sum2[363]==0)Sum2_hex=363;
        else if(Sum2[362]==0)Sum2_hex=362;
        else if(Sum2[361]==0)Sum2_hex=361;
        else if(Sum2[360]==0)Sum2_hex=360;
        else if(Sum2[359]==0)Sum2_hex=359;
        else if(Sum2[358]==0)Sum2_hex=358;
        else if(Sum2[357]==0)Sum2_hex=357;
        else if(Sum2[356]==0)Sum2_hex=356;
        else if(Sum2[355]==0)Sum2_hex=355;
        else if(Sum2[354]==0)Sum2_hex=354;
        else if(Sum2[353]==0)Sum2_hex=353;
        else if(Sum2[352]==0)Sum2_hex=352;
        else if(Sum2[351]==0)Sum2_hex=351;
        else if(Sum2[350]==0)Sum2_hex=350;
        else if(Sum2[349]==0)Sum2_hex=349;
        else if(Sum2[348]==0)Sum2_hex=348;
        else if(Sum2[347]==0)Sum2_hex=347;
        else if(Sum2[346]==0)Sum2_hex=346;
        else if(Sum2[345]==0)Sum2_hex=345;
        else if(Sum2[344]==0)Sum2_hex=344;
        else if(Sum2[343]==0)Sum2_hex=343;
        else if(Sum2[342]==0)Sum2_hex=342;
        else if(Sum2[341]==0)Sum2_hex=341;
        else if(Sum2[340]==0)Sum2_hex=340;
        else if(Sum2[339]==0)Sum2_hex=339;
        else if(Sum2[338]==0)Sum2_hex=338;
        else if(Sum2[337]==0)Sum2_hex=337;
        else if(Sum2[336]==0)Sum2_hex=336;
        else if(Sum2[335]==0)Sum2_hex=335;
        else if(Sum2[334]==0)Sum2_hex=334;
        else if(Sum2[333]==0)Sum2_hex=333;
        else if(Sum2[332]==0)Sum2_hex=332;
        else if(Sum2[331]==0)Sum2_hex=331;
        else if(Sum2[330]==0)Sum2_hex=330;
        else if(Sum2[329]==0)Sum2_hex=329;
        else if(Sum2[328]==0)Sum2_hex=328;
        else if(Sum2[327]==0)Sum2_hex=327;
        else if(Sum2[326]==0)Sum2_hex=326;
        else if(Sum2[325]==0)Sum2_hex=325;
        else if(Sum2[324]==0)Sum2_hex=324;
        else if(Sum2[323]==0)Sum2_hex=323;
        else if(Sum2[322]==0)Sum2_hex=322;
        else if(Sum2[321]==0)Sum2_hex=321;
        else if(Sum2[320]==0)Sum2_hex=320;
        else if(Sum2[319]==0)Sum2_hex=319;
        else if(Sum2[318]==0)Sum2_hex=318;
        else if(Sum2[317]==0)Sum2_hex=317;
        else if(Sum2[316]==0)Sum2_hex=316;
        else if(Sum2[315]==0)Sum2_hex=315;
        else if(Sum2[314]==0)Sum2_hex=314;
        else if(Sum2[313]==0)Sum2_hex=313;
        else if(Sum2[312]==0)Sum2_hex=312;
        else if(Sum2[311]==0)Sum2_hex=311;
        else if(Sum2[310]==0)Sum2_hex=310;
        else if(Sum2[309]==0)Sum2_hex=309;
        else if(Sum2[308]==0)Sum2_hex=308;
        else if(Sum2[307]==0)Sum2_hex=307;
        else if(Sum2[306]==0)Sum2_hex=306;
        else if(Sum2[305]==0)Sum2_hex=305;
        else if(Sum2[304]==0)Sum2_hex=304;
        else if(Sum2[303]==0)Sum2_hex=303;
        else if(Sum2[302]==0)Sum2_hex=302;
        else if(Sum2[301]==0)Sum2_hex=301;
        else if(Sum2[300]==0)Sum2_hex=300;
        else if(Sum2[299]==0)Sum2_hex=299;
        else if(Sum2[298]==0)Sum2_hex=298;
        else if(Sum2[297]==0)Sum2_hex=297;
        else if(Sum2[296]==0)Sum2_hex=296;
        else if(Sum2[295]==0)Sum2_hex=295;
        else if(Sum2[294]==0)Sum2_hex=294;
        else if(Sum2[293]==0)Sum2_hex=293;
        else if(Sum2[292]==0)Sum2_hex=292;
        else if(Sum2[291]==0)Sum2_hex=291;
        else if(Sum2[290]==0)Sum2_hex=290;
        else if(Sum2[289]==0)Sum2_hex=289;
        else if(Sum2[288]==0)Sum2_hex=288;
        else if(Sum2[287]==0)Sum2_hex=287;
        else if(Sum2[286]==0)Sum2_hex=286;
        else if(Sum2[285]==0)Sum2_hex=285;
        else if(Sum2[284]==0)Sum2_hex=284;
        else if(Sum2[283]==0)Sum2_hex=283;
        else if(Sum2[282]==0)Sum2_hex=282;
        else if(Sum2[281]==0)Sum2_hex=281;
        else if(Sum2[280]==0)Sum2_hex=280;
        else if(Sum2[279]==0)Sum2_hex=279;
        else if(Sum2[278]==0)Sum2_hex=278;
        else if(Sum2[277]==0)Sum2_hex=277;
        else if(Sum2[276]==0)Sum2_hex=276;
        else if(Sum2[275]==0)Sum2_hex=275;
        else if(Sum2[274]==0)Sum2_hex=274;
        else if(Sum2[273]==0)Sum2_hex=273;
        else if(Sum2[272]==0)Sum2_hex=272;
        else if(Sum2[271]==0)Sum2_hex=271;
        else if(Sum2[270]==0)Sum2_hex=270;
        else if(Sum2[269]==0)Sum2_hex=269;
        else if(Sum2[268]==0)Sum2_hex=268;
        else if(Sum2[267]==0)Sum2_hex=267;
        else if(Sum2[266]==0)Sum2_hex=266;
        else if(Sum2[265]==0)Sum2_hex=265;
        else if(Sum2[264]==0)Sum2_hex=264;
        else if(Sum2[263]==0)Sum2_hex=263;
        else if(Sum2[262]==0)Sum2_hex=262;
        else if(Sum2[261]==0)Sum2_hex=261;
        else if(Sum2[260]==0)Sum2_hex=260;
        else if(Sum2[259]==0)Sum2_hex=259;
        else if(Sum2[258]==0)Sum2_hex=258;
        else if(Sum2[257]==0)Sum2_hex=257;
        else if(Sum2[256]==0)Sum2_hex=256;
        else if(Sum2[255]==0)Sum2_hex=255;
        else if(Sum2[254]==0)Sum2_hex=254;
        else if(Sum2[253]==0)Sum2_hex=253;
        else if(Sum2[252]==0)Sum2_hex=252;
        else if(Sum2[251]==0)Sum2_hex=251;
        else if(Sum2[250]==0)Sum2_hex=250;
        else if(Sum2[249]==0)Sum2_hex=249;
        else if(Sum2[248]==0)Sum2_hex=248;
        else if(Sum2[247]==0)Sum2_hex=247;
        else if(Sum2[246]==0)Sum2_hex=246;
        else if(Sum2[245]==0)Sum2_hex=245;
        else if(Sum2[244]==0)Sum2_hex=244;
        else if(Sum2[243]==0)Sum2_hex=243;
        else if(Sum2[242]==0)Sum2_hex=242;
        else if(Sum2[241]==0)Sum2_hex=241;
        else if(Sum2[240]==0)Sum2_hex=240;
        else if(Sum2[239]==0)Sum2_hex=239;
        else if(Sum2[238]==0)Sum2_hex=238;
        else if(Sum2[237]==0)Sum2_hex=237;
        else if(Sum2[236]==0)Sum2_hex=236;
        else if(Sum2[235]==0)Sum2_hex=235;
        else if(Sum2[234]==0)Sum2_hex=234;
        else if(Sum2[233]==0)Sum2_hex=233;
        else if(Sum2[232]==0)Sum2_hex=232;
        else if(Sum2[231]==0)Sum2_hex=231;
        else if(Sum2[230]==0)Sum2_hex=230;
        else if(Sum2[229]==0)Sum2_hex=229;
        else if(Sum2[228]==0)Sum2_hex=228;
        else if(Sum2[227]==0)Sum2_hex=227;
        else if(Sum2[226]==0)Sum2_hex=226;
        else if(Sum2[225]==0)Sum2_hex=225;
        else if(Sum2[224]==0)Sum2_hex=224;
        else if(Sum2[223]==0)Sum2_hex=223;
        else if(Sum2[222]==0)Sum2_hex=222;
        else if(Sum2[221]==0)Sum2_hex=221;
        else if(Sum2[220]==0)Sum2_hex=220;
        else if(Sum2[219]==0)Sum2_hex=219;
        else if(Sum2[218]==0)Sum2_hex=218;
        else if(Sum2[217]==0)Sum2_hex=217;
        else if(Sum2[216]==0)Sum2_hex=216;
        else if(Sum2[215]==0)Sum2_hex=215;
        else if(Sum2[214]==0)Sum2_hex=214;
        else if(Sum2[213]==0)Sum2_hex=213;
        else if(Sum2[212]==0)Sum2_hex=212;
        else if(Sum2[211]==0)Sum2_hex=211;
        else if(Sum2[210]==0)Sum2_hex=210;
        else if(Sum2[209]==0)Sum2_hex=209;
        else if(Sum2[208]==0)Sum2_hex=208;
        else if(Sum2[207]==0)Sum2_hex=207;
        else if(Sum2[206]==0)Sum2_hex=206;
        else if(Sum2[205]==0)Sum2_hex=205;
        else if(Sum2[204]==0)Sum2_hex=204;
        else if(Sum2[203]==0)Sum2_hex=203;
        else if(Sum2[202]==0)Sum2_hex=202;
        else if(Sum2[201]==0)Sum2_hex=201;
        else if(Sum2[200]==0)Sum2_hex=200;
        else if(Sum2[199]==0)Sum2_hex=199;
        else if(Sum2[198]==0)Sum2_hex=198;
        else if(Sum2[197]==0)Sum2_hex=197;
        else if(Sum2[196]==0)Sum2_hex=196;
        else if(Sum2[195]==0)Sum2_hex=195;
        else if(Sum2[194]==0)Sum2_hex=194;
        else if(Sum2[193]==0)Sum2_hex=193;
        else if(Sum2[192]==0)Sum2_hex=192;
        else if(Sum2[191]==0)Sum2_hex=191;
        else if(Sum2[190]==0)Sum2_hex=190;
        else if(Sum2[189]==0)Sum2_hex=189;
        else if(Sum2[188]==0)Sum2_hex=188;
        else if(Sum2[187]==0)Sum2_hex=187;
        else if(Sum2[186]==0)Sum2_hex=186;
        else if(Sum2[185]==0)Sum2_hex=185;
        else if(Sum2[184]==0)Sum2_hex=184;
        else if(Sum2[183]==0)Sum2_hex=183;
        else if(Sum2[182]==0)Sum2_hex=182;
        else if(Sum2[181]==0)Sum2_hex=181;
        else if(Sum2[180]==0)Sum2_hex=180;
        else if(Sum2[179]==0)Sum2_hex=179;
        else if(Sum2[178]==0)Sum2_hex=178;
        else if(Sum2[177]==0)Sum2_hex=177;
        else if(Sum2[176]==0)Sum2_hex=176;
        else if(Sum2[175]==0)Sum2_hex=175;
        else if(Sum2[174]==0)Sum2_hex=174;
        else if(Sum2[173]==0)Sum2_hex=173;
        else if(Sum2[172]==0)Sum2_hex=172;
        else if(Sum2[171]==0)Sum2_hex=171;
        else if(Sum2[170]==0)Sum2_hex=170;
        else if(Sum2[169]==0)Sum2_hex=169;
        else if(Sum2[168]==0)Sum2_hex=168;
        else if(Sum2[167]==0)Sum2_hex=167;
        else if(Sum2[166]==0)Sum2_hex=166;
        else if(Sum2[165]==0)Sum2_hex=165;
        else if(Sum2[164]==0)Sum2_hex=164;
        else if(Sum2[163]==0)Sum2_hex=163;
        else if(Sum2[162]==0)Sum2_hex=162;
        else if(Sum2[161]==0)Sum2_hex=161;
        else if(Sum2[160]==0)Sum2_hex=160;
        else if(Sum2[159]==0)Sum2_hex=159;
        else if(Sum2[158]==0)Sum2_hex=158;
        else if(Sum2[157]==0)Sum2_hex=157;
        else if(Sum2[156]==0)Sum2_hex=156;
        else if(Sum2[155]==0)Sum2_hex=155;
        else if(Sum2[154]==0)Sum2_hex=154;
        else if(Sum2[153]==0)Sum2_hex=153;
        else if(Sum2[152]==0)Sum2_hex=152;
        else if(Sum2[151]==0)Sum2_hex=151;
        else if(Sum2[150]==0)Sum2_hex=150;
        else if(Sum2[149]==0)Sum2_hex=149;
        else if(Sum2[148]==0)Sum2_hex=148;
        else if(Sum2[147]==0)Sum2_hex=147;
        else if(Sum2[146]==0)Sum2_hex=146;
        else if(Sum2[145]==0)Sum2_hex=145;
        else if(Sum2[144]==0)Sum2_hex=144;
        else if(Sum2[143]==0)Sum2_hex=143;
        else if(Sum2[142]==0)Sum2_hex=142;
        else if(Sum2[141]==0)Sum2_hex=141;
        else if(Sum2[140]==0)Sum2_hex=140;
        else if(Sum2[139]==0)Sum2_hex=139;
        else if(Sum2[138]==0)Sum2_hex=138;
        else if(Sum2[137]==0)Sum2_hex=137;
        else if(Sum2[136]==0)Sum2_hex=136;
        else if(Sum2[135]==0)Sum2_hex=135;
        else if(Sum2[134]==0)Sum2_hex=134;
        else if(Sum2[133]==0)Sum2_hex=133;
        else if(Sum2[132]==0)Sum2_hex=132;
        else if(Sum2[131]==0)Sum2_hex=131;
        else if(Sum2[130]==0)Sum2_hex=130;
        else if(Sum2[129]==0)Sum2_hex=129;
        else if(Sum2[128]==0)Sum2_hex=128;
        else if(Sum2[127]==0)Sum2_hex=127;
        else if(Sum2[126]==0)Sum2_hex=126;
        else if(Sum2[125]==0)Sum2_hex=125;
        else if(Sum2[124]==0)Sum2_hex=124;
        else if(Sum2[123]==0)Sum2_hex=123;
        else if(Sum2[122]==0)Sum2_hex=122;
        else if(Sum2[121]==0)Sum2_hex=121;
        else if(Sum2[120]==0)Sum2_hex=120;
        else if(Sum2[119]==0)Sum2_hex=119;
        else if(Sum2[118]==0)Sum2_hex=118;
        else if(Sum2[117]==0)Sum2_hex=117;
        else if(Sum2[116]==0)Sum2_hex=116;
        else if(Sum2[115]==0)Sum2_hex=115;
        else if(Sum2[114]==0)Sum2_hex=114;
        else if(Sum2[113]==0)Sum2_hex=113;
        else if(Sum2[112]==0)Sum2_hex=112;
        else if(Sum2[111]==0)Sum2_hex=111;
        else if(Sum2[110]==0)Sum2_hex=110;
        else if(Sum2[109]==0)Sum2_hex=109;
        else if(Sum2[108]==0)Sum2_hex=108;
        else if(Sum2[107]==0)Sum2_hex=107;
        else if(Sum2[106]==0)Sum2_hex=106;
        else if(Sum2[105]==0)Sum2_hex=105;
        else if(Sum2[104]==0)Sum2_hex=104;
        else if(Sum2[103]==0)Sum2_hex=103;
        else if(Sum2[102]==0)Sum2_hex=102;
        else if(Sum2[101]==0)Sum2_hex=101;
        else if(Sum2[100]==0)Sum2_hex=100;
        else if(Sum2[99]==0)Sum2_hex=99;
        else if(Sum2[98]==0)Sum2_hex=98;
        else if(Sum2[97]==0)Sum2_hex=97;
        else if(Sum2[96]==0)Sum2_hex=96;
        else if(Sum2[95]==0)Sum2_hex=95;
        else if(Sum2[94]==0)Sum2_hex=94;
        else if(Sum2[93]==0)Sum2_hex=93;
        else if(Sum2[92]==0)Sum2_hex=92;
        else if(Sum2[91]==0)Sum2_hex=91;
        else if(Sum2[90]==0)Sum2_hex=90;
        else if(Sum2[89]==0)Sum2_hex=89;
        else if(Sum2[88]==0)Sum2_hex=88;
        else if(Sum2[87]==0)Sum2_hex=87;
        else if(Sum2[86]==0)Sum2_hex=86;
        else if(Sum2[85]==0)Sum2_hex=85;
        else if(Sum2[84]==0)Sum2_hex=84;
        else if(Sum2[83]==0)Sum2_hex=83;
        else if(Sum2[82]==0)Sum2_hex=82;
        else if(Sum2[81]==0)Sum2_hex=81;
        else if(Sum2[80]==0)Sum2_hex=80;
        else if(Sum2[79]==0)Sum2_hex=79;
        else if(Sum2[78]==0)Sum2_hex=78;
        else if(Sum2[77]==0)Sum2_hex=77;
        else if(Sum2[76]==0)Sum2_hex=76;
        else if(Sum2[75]==0)Sum2_hex=75;
        else if(Sum2[74]==0)Sum2_hex=74;
        else if(Sum2[73]==0)Sum2_hex=73;
        else if(Sum2[72]==0)Sum2_hex=72;
        else if(Sum2[71]==0)Sum2_hex=71;
        else if(Sum2[70]==0)Sum2_hex=70;
        else if(Sum2[69]==0)Sum2_hex=69;
        else if(Sum2[68]==0)Sum2_hex=68;
        else if(Sum2[67]==0)Sum2_hex=67;
        else if(Sum2[66]==0)Sum2_hex=66;
        else if(Sum2[65]==0)Sum2_hex=65;
        else if(Sum2[64]==0)Sum2_hex=64;
        else if(Sum2[63]==0)Sum2_hex=63;
        else if(Sum2[62]==0)Sum2_hex=62;
        else if(Sum2[61]==0)Sum2_hex=61;
        else if(Sum2[60]==0)Sum2_hex=60;
        else if(Sum2[59]==0)Sum2_hex=59;
        else if(Sum2[58]==0)Sum2_hex=58;
        else if(Sum2[57]==0)Sum2_hex=57;
        else if(Sum2[56]==0)Sum2_hex=56;
        else if(Sum2[55]==0)Sum2_hex=55;
        else if(Sum2[54]==0)Sum2_hex=54;
        else if(Sum2[53]==0)Sum2_hex=53;
        else if(Sum2[52]==0)Sum2_hex=52;
        else if(Sum2[51]==0)Sum2_hex=51;
        else if(Sum2[50]==0)Sum2_hex=50;
        else if(Sum2[49]==0)Sum2_hex=49;
        else if(Sum2[48]==0)Sum2_hex=48;
        else if(Sum2[47]==0)Sum2_hex=47;
        else if(Sum2[46]==0)Sum2_hex=46;
        else if(Sum2[45]==0)Sum2_hex=45;
        else if(Sum2[44]==0)Sum2_hex=44;
        else if(Sum2[43]==0)Sum2_hex=43;
        else if(Sum2[42]==0)Sum2_hex=42;
        else if(Sum2[41]==0)Sum2_hex=41;
        else if(Sum2[40]==0)Sum2_hex=40;
        else if(Sum2[39]==0)Sum2_hex=39;
        else if(Sum2[38]==0)Sum2_hex=38;
        else if(Sum2[37]==0)Sum2_hex=37;
        else if(Sum2[36]==0)Sum2_hex=36;
        else if(Sum2[35]==0)Sum2_hex=35;
        else if(Sum2[34]==0)Sum2_hex=34;
        else if(Sum2[33]==0)Sum2_hex=33;
        else if(Sum2[32]==0)Sum2_hex=32;
        else if(Sum2[31]==0)Sum2_hex=31;
        else if(Sum2[30]==0)Sum2_hex=30;
        else if(Sum2[29]==0)Sum2_hex=29;
        else if(Sum2[28]==0)Sum2_hex=28;
        else if(Sum2[27]==0)Sum2_hex=27;
        else if(Sum2[26]==0)Sum2_hex=26;
        else if(Sum2[25]==0)Sum2_hex=25;
        else if(Sum2[24]==0)Sum2_hex=24;
        else if(Sum2[23]==0)Sum2_hex=23;
        else if(Sum2[22]==0)Sum2_hex=22;
        else if(Sum2[21]==0)Sum2_hex=21;
        else if(Sum2[20]==0)Sum2_hex=20;
        else if(Sum2[19]==0)Sum2_hex=19;
        else if(Sum2[18]==0)Sum2_hex=18;
        else if(Sum2[17]==0)Sum2_hex=17;
        else if(Sum2[16]==0)Sum2_hex=16;
        else if(Sum2[15]==0)Sum2_hex=15;
        else if(Sum2[14]==0)Sum2_hex=14;
        else if(Sum2[13]==0)Sum2_hex=13;
        else if(Sum2[12]==0)Sum2_hex=12;
        else if(Sum2[11]==0)Sum2_hex=11;
        else if(Sum2[10]==0)Sum2_hex=10;
        else if(Sum2[9]==0)Sum2_hex=9;
        else if(Sum2[8]==0)Sum2_hex=8;
        else if(Sum2[7]==0)Sum2_hex=7;
        else if(Sum2[6]==0)Sum2_hex=6;
        else if(Sum2[5]==0)Sum2_hex=5;
        else if(Sum2[4]==0)Sum2_hex=4;
        else if(Sum2[3]==0)Sum2_hex=3;
        else if(Sum2[2]==0)Sum2_hex=2;
        else if(Sum2[1]==0)Sum2_hex=1;
        else if(Sum2[0]==0)Sum2_hex=0;
        else Sum2_hex=0;
    end
    else begin
        Sum2_hex=2184;
    end
end

always @(posedge Hit) begin 
        Sum2[1023:0] <= 4096'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
        Co2[1023:0] <= 4096'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        Sum2[0]<=1^Hit^Ci;
        Co2[0]<=(1&Hit|(1|Hit)&Ci);

        Sum2[1]<=1^0^Co2[0];
        Co2[1]<=(1&0|(1|0)&Co2[0]);

        Sum2[2]<=1^0^Co2[1];
        Co2[2]<=(1&0|(1|0)&Co2[1]);

        Sum2[3]<=1^0^Co2[2];
        Co2[3]<=(1&0|(1|0)&Co2[2]);

        Sum2[4]<=1^0^Co2[3];
        Co2[4]<=(1&0|(1|0)&Co2[3]);

        Sum2[5]<=1^0^Co2[4];
        Co2[5]<=(1&0|(1|0)&Co2[4]);

        Sum2[6]<=1^0^Co2[5];
        Co2[6]<=(1&0|(1|0)&Co2[5]);

        Sum2[7]<=1^0^Co2[6];
        Co2[7]<=(1&0|(1|0)&Co2[6]);

        Sum2[8]<=1^0^Co2[7];
        Co2[8]<=(1&0|(1|0)&Co2[7]);

        Sum2[9]<=1^0^Co2[8];
        Co2[9]<=(1&0|(1|0)&Co2[8]);

        Sum2[10]<=1^0^Co2[9];
        Co2[10]<=(1&0|(1|0)&Co2[9]);

        Sum2[11]<=1^0^Co2[10];
        Co2[11]<=(1&0|(1|0)&Co2[10]);

        Sum2[12]<=1^0^Co2[11];
        Co2[12]<=(1&0|(1|0)&Co2[11]);

        Sum2[13]<=1^0^Co2[12];
        Co2[13]<=(1&0|(1|0)&Co2[12]);

        Sum2[14]<=1^0^Co2[13];
        Co2[14]<=(1&0|(1|0)&Co2[13]);

        Sum2[15]<=1^0^Co2[14];
        Co2[15]<=(1&0|(1|0)&Co2[14]);

        Sum2[16]<=1^0^Co2[15];
        Co2[16]<=(1&0|(1|0)&Co2[15]);

        Sum2[17]<=1^0^Co2[16];
        Co2[17]<=(1&0|(1|0)&Co2[16]);

        Sum2[18]<=1^0^Co2[17];
        Co2[18]<=(1&0|(1|0)&Co2[17]);

        Sum2[19]<=1^0^Co2[18];
        Co2[19]<=(1&0|(1|0)&Co2[18]);

        Sum2[20]<=1^0^Co2[19];
        Co2[20]<=(1&0|(1|0)&Co2[19]);

        Sum2[21]<=1^0^Co2[20];
        Co2[21]<=(1&0|(1|0)&Co2[20]);

        Sum2[22]<=1^0^Co2[21];
        Co2[22]<=(1&0|(1|0)&Co2[21]);

        Sum2[23]<=1^0^Co2[22];
        Co2[23]<=(1&0|(1|0)&Co2[22]);

        Sum2[24]<=1^0^Co2[23];
        Co2[24]<=(1&0|(1|0)&Co2[23]);

        Sum2[25]<=1^0^Co2[24];
        Co2[25]<=(1&0|(1|0)&Co2[24]);

        Sum2[26]<=1^0^Co2[25];
        Co2[26]<=(1&0|(1|0)&Co2[25]);

        Sum2[27]<=1^0^Co2[26];
        Co2[27]<=(1&0|(1|0)&Co2[26]);

        Sum2[28]<=1^0^Co2[27];
        Co2[28]<=(1&0|(1|0)&Co2[27]);

        Sum2[29]<=1^0^Co2[28];
        Co2[29]<=(1&0|(1|0)&Co2[28]);

        Sum2[30]<=1^0^Co2[29];
        Co2[30]<=(1&0|(1|0)&Co2[29]);

        Sum2[31]<=1^0^Co2[30];
        Co2[31]<=(1&0|(1|0)&Co2[30]);

        Sum2[32]<=1^0^Co2[31];
        Co2[32]<=(1&0|(1|0)&Co2[31]);

        Sum2[33]<=1^0^Co2[32];
        Co2[33]<=(1&0|(1|0)&Co2[32]);

        Sum2[34]<=1^0^Co2[33];
        Co2[34]<=(1&0|(1|0)&Co2[33]);

        Sum2[35]<=1^0^Co2[34];
        Co2[35]<=(1&0|(1|0)&Co2[34]);

        Sum2[36]<=1^0^Co2[35];
        Co2[36]<=(1&0|(1|0)&Co2[35]);

        Sum2[37]<=1^0^Co2[36];
        Co2[37]<=(1&0|(1|0)&Co2[36]);

        Sum2[38]<=1^0^Co2[37];
        Co2[38]<=(1&0|(1|0)&Co2[37]);

        Sum2[39]<=1^0^Co2[38];
        Co2[39]<=(1&0|(1|0)&Co2[38]);

        Sum2[40]<=1^0^Co2[39];
        Co2[40]<=(1&0|(1|0)&Co2[39]);

        Sum2[41]<=1^0^Co2[40];
        Co2[41]<=(1&0|(1|0)&Co2[40]);

        Sum2[42]<=1^0^Co2[41];
        Co2[42]<=(1&0|(1|0)&Co2[41]);

        Sum2[43]<=1^0^Co2[42];
        Co2[43]<=(1&0|(1|0)&Co2[42]);

        Sum2[44]<=1^0^Co2[43];
        Co2[44]<=(1&0|(1|0)&Co2[43]);

        Sum2[45]<=1^0^Co2[44];
        Co2[45]<=(1&0|(1|0)&Co2[44]);

        Sum2[46]<=1^0^Co2[45];
        Co2[46]<=(1&0|(1|0)&Co2[45]);

        Sum2[47]<=1^0^Co2[46];
        Co2[47]<=(1&0|(1|0)&Co2[46]);

        Sum2[48]<=1^0^Co2[47];
        Co2[48]<=(1&0|(1|0)&Co2[47]);

        Sum2[49]<=1^0^Co2[48];
        Co2[49]<=(1&0|(1|0)&Co2[48]);

        Sum2[50]<=1^0^Co2[49];
        Co2[50]<=(1&0|(1|0)&Co2[49]);

        Sum2[51]<=1^0^Co2[50];
        Co2[51]<=(1&0|(1|0)&Co2[50]);

        Sum2[52]<=1^0^Co2[51];
        Co2[52]<=(1&0|(1|0)&Co2[51]);

        Sum2[53]<=1^0^Co2[52];
        Co2[53]<=(1&0|(1|0)&Co2[52]);

        Sum2[54]<=1^0^Co2[53];
        Co2[54]<=(1&0|(1|0)&Co2[53]);

        Sum2[55]<=1^0^Co2[54];
        Co2[55]<=(1&0|(1|0)&Co2[54]);

        Sum2[56]<=1^0^Co2[55];
        Co2[56]<=(1&0|(1|0)&Co2[55]);

        Sum2[57]<=1^0^Co2[56];
        Co2[57]<=(1&0|(1|0)&Co2[56]);

        Sum2[58]<=1^0^Co2[57];
        Co2[58]<=(1&0|(1|0)&Co2[57]);

        Sum2[59]<=1^0^Co2[58];
        Co2[59]<=(1&0|(1|0)&Co2[58]);

        Sum2[60]<=1^0^Co2[59];
        Co2[60]<=(1&0|(1|0)&Co2[59]);

        Sum2[61]<=1^0^Co2[60];
        Co2[61]<=(1&0|(1|0)&Co2[60]);

        Sum2[62]<=1^0^Co2[61];
        Co2[62]<=(1&0|(1|0)&Co2[61]);

        Sum2[63]<=1^0^Co2[62];
        Co2[63]<=(1&0|(1|0)&Co2[62]);

        Sum2[64]<=1^0^Co2[63];
        Co2[64]<=(1&0|(1|0)&Co2[63]);

        Sum2[65]<=1^0^Co2[64];
        Co2[65]<=(1&0|(1|0)&Co2[64]);

        Sum2[66]<=1^0^Co2[65];
        Co2[66]<=(1&0|(1|0)&Co2[65]);

        Sum2[67]<=1^0^Co2[66];
        Co2[67]<=(1&0|(1|0)&Co2[66]);

        Sum2[68]<=1^0^Co2[67];
        Co2[68]<=(1&0|(1|0)&Co2[67]);

        Sum2[69]<=1^0^Co2[68];
        Co2[69]<=(1&0|(1|0)&Co2[68]);

        Sum2[70]<=1^0^Co2[69];
        Co2[70]<=(1&0|(1|0)&Co2[69]);

        Sum2[71]<=1^0^Co2[70];
        Co2[71]<=(1&0|(1|0)&Co2[70]);

        Sum2[72]<=1^0^Co2[71];
        Co2[72]<=(1&0|(1|0)&Co2[71]);

        Sum2[73]<=1^0^Co2[72];
        Co2[73]<=(1&0|(1|0)&Co2[72]);

        Sum2[74]<=1^0^Co2[73];
        Co2[74]<=(1&0|(1|0)&Co2[73]);

        Sum2[75]<=1^0^Co2[74];
        Co2[75]<=(1&0|(1|0)&Co2[74]);

        Sum2[76]<=1^0^Co2[75];
        Co2[76]<=(1&0|(1|0)&Co2[75]);

        Sum2[77]<=1^0^Co2[76];
        Co2[77]<=(1&0|(1|0)&Co2[76]);

        Sum2[78]<=1^0^Co2[77];
        Co2[78]<=(1&0|(1|0)&Co2[77]);

        Sum2[79]<=1^0^Co2[78];
        Co2[79]<=(1&0|(1|0)&Co2[78]);

        Sum2[80]<=1^0^Co2[79];
        Co2[80]<=(1&0|(1|0)&Co2[79]);

        Sum2[81]<=1^0^Co2[80];
        Co2[81]<=(1&0|(1|0)&Co2[80]);

        Sum2[82]<=1^0^Co2[81];
        Co2[82]<=(1&0|(1|0)&Co2[81]);

        Sum2[83]<=1^0^Co2[82];
        Co2[83]<=(1&0|(1|0)&Co2[82]);

        Sum2[84]<=1^0^Co2[83];
        Co2[84]<=(1&0|(1|0)&Co2[83]);

        Sum2[85]<=1^0^Co2[84];
        Co2[85]<=(1&0|(1|0)&Co2[84]);

        Sum2[86]<=1^0^Co2[85];
        Co2[86]<=(1&0|(1|0)&Co2[85]);

        Sum2[87]<=1^0^Co2[86];
        Co2[87]<=(1&0|(1|0)&Co2[86]);

        Sum2[88]<=1^0^Co2[87];
        Co2[88]<=(1&0|(1|0)&Co2[87]);

        Sum2[89]<=1^0^Co2[88];
        Co2[89]<=(1&0|(1|0)&Co2[88]);

        Sum2[90]<=1^0^Co2[89];
        Co2[90]<=(1&0|(1|0)&Co2[89]);

        Sum2[91]<=1^0^Co2[90];
        Co2[91]<=(1&0|(1|0)&Co2[90]);

        Sum2[92]<=1^0^Co2[91];
        Co2[92]<=(1&0|(1|0)&Co2[91]);

        Sum2[93]<=1^0^Co2[92];
        Co2[93]<=(1&0|(1|0)&Co2[92]);

        Sum2[94]<=1^0^Co2[93];
        Co2[94]<=(1&0|(1|0)&Co2[93]);

        Sum2[95]<=1^0^Co2[94];
        Co2[95]<=(1&0|(1|0)&Co2[94]);

        Sum2[96]<=1^0^Co2[95];
        Co2[96]<=(1&0|(1|0)&Co2[95]);

        Sum2[97]<=1^0^Co2[96];
        Co2[97]<=(1&0|(1|0)&Co2[96]);

        Sum2[98]<=1^0^Co2[97];
        Co2[98]<=(1&0|(1|0)&Co2[97]);

        Sum2[99]<=1^0^Co2[98];
        Co2[99]<=(1&0|(1|0)&Co2[98]);

        Sum2[100]<=1^0^Co2[99];
        Co2[100]<=(1&0|(1|0)&Co2[99]);

        Sum2[101]<=1^0^Co2[100];
        Co2[101]<=(1&0|(1|0)&Co2[100]);

        Sum2[102]<=1^0^Co2[101];
        Co2[102]<=(1&0|(1|0)&Co2[101]);

        Sum2[103]<=1^0^Co2[102];
        Co2[103]<=(1&0|(1|0)&Co2[102]);

        Sum2[104]<=1^0^Co2[103];
        Co2[104]<=(1&0|(1|0)&Co2[103]);

        Sum2[105]<=1^0^Co2[104];
        Co2[105]<=(1&0|(1|0)&Co2[104]);

        Sum2[106]<=1^0^Co2[105];
        Co2[106]<=(1&0|(1|0)&Co2[105]);

        Sum2[107]<=1^0^Co2[106];
        Co2[107]<=(1&0|(1|0)&Co2[106]);

        Sum2[108]<=1^0^Co2[107];
        Co2[108]<=(1&0|(1|0)&Co2[107]);

        Sum2[109]<=1^0^Co2[108];
        Co2[109]<=(1&0|(1|0)&Co2[108]);

        Sum2[110]<=1^0^Co2[109];
        Co2[110]<=(1&0|(1|0)&Co2[109]);

        Sum2[111]<=1^0^Co2[110];
        Co2[111]<=(1&0|(1|0)&Co2[110]);

        Sum2[112]<=1^0^Co2[111];
        Co2[112]<=(1&0|(1|0)&Co2[111]);

        Sum2[113]<=1^0^Co2[112];
        Co2[113]<=(1&0|(1|0)&Co2[112]);

        Sum2[114]<=1^0^Co2[113];
        Co2[114]<=(1&0|(1|0)&Co2[113]);

        Sum2[115]<=1^0^Co2[114];
        Co2[115]<=(1&0|(1|0)&Co2[114]);

        Sum2[116]<=1^0^Co2[115];
        Co2[116]<=(1&0|(1|0)&Co2[115]);

        Sum2[117]<=1^0^Co2[116];
        Co2[117]<=(1&0|(1|0)&Co2[116]);

        Sum2[118]<=1^0^Co2[117];
        Co2[118]<=(1&0|(1|0)&Co2[117]);

        Sum2[119]<=1^0^Co2[118];
        Co2[119]<=(1&0|(1|0)&Co2[118]);

        Sum2[120]<=1^0^Co2[119];
        Co2[120]<=(1&0|(1|0)&Co2[119]);

        Sum2[121]<=1^0^Co2[120];
        Co2[121]<=(1&0|(1|0)&Co2[120]);

        Sum2[122]<=1^0^Co2[121];
        Co2[122]<=(1&0|(1|0)&Co2[121]);

        Sum2[123]<=1^0^Co2[122];
        Co2[123]<=(1&0|(1|0)&Co2[122]);

        Sum2[124]<=1^0^Co2[123];
        Co2[124]<=(1&0|(1|0)&Co2[123]);

        Sum2[125]<=1^0^Co2[124];
        Co2[125]<=(1&0|(1|0)&Co2[124]);

        Sum2[126]<=1^0^Co2[125];
        Co2[126]<=(1&0|(1|0)&Co2[125]);

        Sum2[127]<=1^0^Co2[126];
        Co2[127]<=(1&0|(1|0)&Co2[126]);

        Sum2[128]<=1^0^Co2[127];
        Co2[128]<=(1&0|(1|0)&Co2[127]);

        Sum2[129]<=1^0^Co2[128];
        Co2[129]<=(1&0|(1|0)&Co2[128]);

        Sum2[130]<=1^0^Co2[129];
        Co2[130]<=(1&0|(1|0)&Co2[129]);

        Sum2[131]<=1^0^Co2[130];
        Co2[131]<=(1&0|(1|0)&Co2[130]);

        Sum2[132]<=1^0^Co2[131];
        Co2[132]<=(1&0|(1|0)&Co2[131]);

        Sum2[133]<=1^0^Co2[132];
        Co2[133]<=(1&0|(1|0)&Co2[132]);

        Sum2[134]<=1^0^Co2[133];
        Co2[134]<=(1&0|(1|0)&Co2[133]);

        Sum2[135]<=1^0^Co2[134];
        Co2[135]<=(1&0|(1|0)&Co2[134]);

        Sum2[136]<=1^0^Co2[135];
        Co2[136]<=(1&0|(1|0)&Co2[135]);

        Sum2[137]<=1^0^Co2[136];
        Co2[137]<=(1&0|(1|0)&Co2[136]);

        Sum2[138]<=1^0^Co2[137];
        Co2[138]<=(1&0|(1|0)&Co2[137]);

        Sum2[139]<=1^0^Co2[138];
        Co2[139]<=(1&0|(1|0)&Co2[138]);

        Sum2[140]<=1^0^Co2[139];
        Co2[140]<=(1&0|(1|0)&Co2[139]);

        Sum2[141]<=1^0^Co2[140];
        Co2[141]<=(1&0|(1|0)&Co2[140]);

        Sum2[142]<=1^0^Co2[141];
        Co2[142]<=(1&0|(1|0)&Co2[141]);

        Sum2[143]<=1^0^Co2[142];
        Co2[143]<=(1&0|(1|0)&Co2[142]);

        Sum2[144]<=1^0^Co2[143];
        Co2[144]<=(1&0|(1|0)&Co2[143]);

        Sum2[145]<=1^0^Co2[144];
        Co2[145]<=(1&0|(1|0)&Co2[144]);

        Sum2[146]<=1^0^Co2[145];
        Co2[146]<=(1&0|(1|0)&Co2[145]);

        Sum2[147]<=1^0^Co2[146];
        Co2[147]<=(1&0|(1|0)&Co2[146]);

        Sum2[148]<=1^0^Co2[147];
        Co2[148]<=(1&0|(1|0)&Co2[147]);

        Sum2[149]<=1^0^Co2[148];
        Co2[149]<=(1&0|(1|0)&Co2[148]);

        Sum2[150]<=1^0^Co2[149];
        Co2[150]<=(1&0|(1|0)&Co2[149]);

        Sum2[151]<=1^0^Co2[150];
        Co2[151]<=(1&0|(1|0)&Co2[150]);

        Sum2[152]<=1^0^Co2[151];
        Co2[152]<=(1&0|(1|0)&Co2[151]);

        Sum2[153]<=1^0^Co2[152];
        Co2[153]<=(1&0|(1|0)&Co2[152]);

        Sum2[154]<=1^0^Co2[153];
        Co2[154]<=(1&0|(1|0)&Co2[153]);

        Sum2[155]<=1^0^Co2[154];
        Co2[155]<=(1&0|(1|0)&Co2[154]);

        Sum2[156]<=1^0^Co2[155];
        Co2[156]<=(1&0|(1|0)&Co2[155]);

        Sum2[157]<=1^0^Co2[156];
        Co2[157]<=(1&0|(1|0)&Co2[156]);

        Sum2[158]<=1^0^Co2[157];
        Co2[158]<=(1&0|(1|0)&Co2[157]);

        Sum2[159]<=1^0^Co2[158];
        Co2[159]<=(1&0|(1|0)&Co2[158]);

        Sum2[160]<=1^0^Co2[159];
        Co2[160]<=(1&0|(1|0)&Co2[159]);

        Sum2[161]<=1^0^Co2[160];
        Co2[161]<=(1&0|(1|0)&Co2[160]);

        Sum2[162]<=1^0^Co2[161];
        Co2[162]<=(1&0|(1|0)&Co2[161]);

        Sum2[163]<=1^0^Co2[162];
        Co2[163]<=(1&0|(1|0)&Co2[162]);

        Sum2[164]<=1^0^Co2[163];
        Co2[164]<=(1&0|(1|0)&Co2[163]);

        Sum2[165]<=1^0^Co2[164];
        Co2[165]<=(1&0|(1|0)&Co2[164]);

        Sum2[166]<=1^0^Co2[165];
        Co2[166]<=(1&0|(1|0)&Co2[165]);

        Sum2[167]<=1^0^Co2[166];
        Co2[167]<=(1&0|(1|0)&Co2[166]);

        Sum2[168]<=1^0^Co2[167];
        Co2[168]<=(1&0|(1|0)&Co2[167]);

        Sum2[169]<=1^0^Co2[168];
        Co2[169]<=(1&0|(1|0)&Co2[168]);

        Sum2[170]<=1^0^Co2[169];
        Co2[170]<=(1&0|(1|0)&Co2[169]);

        Sum2[171]<=1^0^Co2[170];
        Co2[171]<=(1&0|(1|0)&Co2[170]);

        Sum2[172]<=1^0^Co2[171];
        Co2[172]<=(1&0|(1|0)&Co2[171]);

        Sum2[173]<=1^0^Co2[172];
        Co2[173]<=(1&0|(1|0)&Co2[172]);

        Sum2[174]<=1^0^Co2[173];
        Co2[174]<=(1&0|(1|0)&Co2[173]);

        Sum2[175]<=1^0^Co2[174];
        Co2[175]<=(1&0|(1|0)&Co2[174]);

        Sum2[176]<=1^0^Co2[175];
        Co2[176]<=(1&0|(1|0)&Co2[175]);

        Sum2[177]<=1^0^Co2[176];
        Co2[177]<=(1&0|(1|0)&Co2[176]);

        Sum2[178]<=1^0^Co2[177];
        Co2[178]<=(1&0|(1|0)&Co2[177]);

        Sum2[179]<=1^0^Co2[178];
        Co2[179]<=(1&0|(1|0)&Co2[178]);

        Sum2[180]<=1^0^Co2[179];
        Co2[180]<=(1&0|(1|0)&Co2[179]);

        Sum2[181]<=1^0^Co2[180];
        Co2[181]<=(1&0|(1|0)&Co2[180]);

        Sum2[182]<=1^0^Co2[181];
        Co2[182]<=(1&0|(1|0)&Co2[181]);

        Sum2[183]<=1^0^Co2[182];
        Co2[183]<=(1&0|(1|0)&Co2[182]);

        Sum2[184]<=1^0^Co2[183];
        Co2[184]<=(1&0|(1|0)&Co2[183]);

        Sum2[185]<=1^0^Co2[184];
        Co2[185]<=(1&0|(1|0)&Co2[184]);

        Sum2[186]<=1^0^Co2[185];
        Co2[186]<=(1&0|(1|0)&Co2[185]);

        Sum2[187]<=1^0^Co2[186];
        Co2[187]<=(1&0|(1|0)&Co2[186]);

        Sum2[188]<=1^0^Co2[187];
        Co2[188]<=(1&0|(1|0)&Co2[187]);

        Sum2[189]<=1^0^Co2[188];
        Co2[189]<=(1&0|(1|0)&Co2[188]);

        Sum2[190]<=1^0^Co2[189];
        Co2[190]<=(1&0|(1|0)&Co2[189]);

        Sum2[191]<=1^0^Co2[190];
        Co2[191]<=(1&0|(1|0)&Co2[190]);

        Sum2[192]<=1^0^Co2[191];
        Co2[192]<=(1&0|(1|0)&Co2[191]);

        Sum2[193]<=1^0^Co2[192];
        Co2[193]<=(1&0|(1|0)&Co2[192]);

        Sum2[194]<=1^0^Co2[193];
        Co2[194]<=(1&0|(1|0)&Co2[193]);

        Sum2[195]<=1^0^Co2[194];
        Co2[195]<=(1&0|(1|0)&Co2[194]);

        Sum2[196]<=1^0^Co2[195];
        Co2[196]<=(1&0|(1|0)&Co2[195]);

        Sum2[197]<=1^0^Co2[196];
        Co2[197]<=(1&0|(1|0)&Co2[196]);

        Sum2[198]<=1^0^Co2[197];
        Co2[198]<=(1&0|(1|0)&Co2[197]);

        Sum2[199]<=1^0^Co2[198];
        Co2[199]<=(1&0|(1|0)&Co2[198]);

        Sum2[200]<=1^0^Co2[199];
        Co2[200]<=(1&0|(1|0)&Co2[199]);

        Sum2[201]<=1^0^Co2[200];
        Co2[201]<=(1&0|(1|0)&Co2[200]);

        Sum2[202]<=1^0^Co2[201];
        Co2[202]<=(1&0|(1|0)&Co2[201]);

        Sum2[203]<=1^0^Co2[202];
        Co2[203]<=(1&0|(1|0)&Co2[202]);

        Sum2[204]<=1^0^Co2[203];
        Co2[204]<=(1&0|(1|0)&Co2[203]);

        Sum2[205]<=1^0^Co2[204];
        Co2[205]<=(1&0|(1|0)&Co2[204]);

        Sum2[206]<=1^0^Co2[205];
        Co2[206]<=(1&0|(1|0)&Co2[205]);

        Sum2[207]<=1^0^Co2[206];
        Co2[207]<=(1&0|(1|0)&Co2[206]);

        Sum2[208]<=1^0^Co2[207];
        Co2[208]<=(1&0|(1|0)&Co2[207]);

        Sum2[209]<=1^0^Co2[208];
        Co2[209]<=(1&0|(1|0)&Co2[208]);

        Sum2[210]<=1^0^Co2[209];
        Co2[210]<=(1&0|(1|0)&Co2[209]);

        Sum2[211]<=1^0^Co2[210];
        Co2[211]<=(1&0|(1|0)&Co2[210]);

        Sum2[212]<=1^0^Co2[211];
        Co2[212]<=(1&0|(1|0)&Co2[211]);

        Sum2[213]<=1^0^Co2[212];
        Co2[213]<=(1&0|(1|0)&Co2[212]);

        Sum2[214]<=1^0^Co2[213];
        Co2[214]<=(1&0|(1|0)&Co2[213]);

        Sum2[215]<=1^0^Co2[214];
        Co2[215]<=(1&0|(1|0)&Co2[214]);

        Sum2[216]<=1^0^Co2[215];
        Co2[216]<=(1&0|(1|0)&Co2[215]);

        Sum2[217]<=1^0^Co2[216];
        Co2[217]<=(1&0|(1|0)&Co2[216]);

        Sum2[218]<=1^0^Co2[217];
        Co2[218]<=(1&0|(1|0)&Co2[217]);

        Sum2[219]<=1^0^Co2[218];
        Co2[219]<=(1&0|(1|0)&Co2[218]);

        Sum2[220]<=1^0^Co2[219];
        Co2[220]<=(1&0|(1|0)&Co2[219]);

        Sum2[221]<=1^0^Co2[220];
        Co2[221]<=(1&0|(1|0)&Co2[220]);

        Sum2[222]<=1^0^Co2[221];
        Co2[222]<=(1&0|(1|0)&Co2[221]);

        Sum2[223]<=1^0^Co2[222];
        Co2[223]<=(1&0|(1|0)&Co2[222]);

        Sum2[224]<=1^0^Co2[223];
        Co2[224]<=(1&0|(1|0)&Co2[223]);

        Sum2[225]<=1^0^Co2[224];
        Co2[225]<=(1&0|(1|0)&Co2[224]);

        Sum2[226]<=1^0^Co2[225];
        Co2[226]<=(1&0|(1|0)&Co2[225]);

        Sum2[227]<=1^0^Co2[226];
        Co2[227]<=(1&0|(1|0)&Co2[226]);

        Sum2[228]<=1^0^Co2[227];
        Co2[228]<=(1&0|(1|0)&Co2[227]);

        Sum2[229]<=1^0^Co2[228];
        Co2[229]<=(1&0|(1|0)&Co2[228]);

        Sum2[230]<=1^0^Co2[229];
        Co2[230]<=(1&0|(1|0)&Co2[229]);

        Sum2[231]<=1^0^Co2[230];
        Co2[231]<=(1&0|(1|0)&Co2[230]);

        Sum2[232]<=1^0^Co2[231];
        Co2[232]<=(1&0|(1|0)&Co2[231]);

        Sum2[233]<=1^0^Co2[232];
        Co2[233]<=(1&0|(1|0)&Co2[232]);

        Sum2[234]<=1^0^Co2[233];
        Co2[234]<=(1&0|(1|0)&Co2[233]);

        Sum2[235]<=1^0^Co2[234];
        Co2[235]<=(1&0|(1|0)&Co2[234]);

        Sum2[236]<=1^0^Co2[235];
        Co2[236]<=(1&0|(1|0)&Co2[235]);

        Sum2[237]<=1^0^Co2[236];
        Co2[237]<=(1&0|(1|0)&Co2[236]);

        Sum2[238]<=1^0^Co2[237];
        Co2[238]<=(1&0|(1|0)&Co2[237]);

        Sum2[239]<=1^0^Co2[238];
        Co2[239]<=(1&0|(1|0)&Co2[238]);

        Sum2[240]<=1^0^Co2[239];
        Co2[240]<=(1&0|(1|0)&Co2[239]);

        Sum2[241]<=1^0^Co2[240];
        Co2[241]<=(1&0|(1|0)&Co2[240]);

        Sum2[242]<=1^0^Co2[241];
        Co2[242]<=(1&0|(1|0)&Co2[241]);

        Sum2[243]<=1^0^Co2[242];
        Co2[243]<=(1&0|(1|0)&Co2[242]);

        Sum2[244]<=1^0^Co2[243];
        Co2[244]<=(1&0|(1|0)&Co2[243]);

        Sum2[245]<=1^0^Co2[244];
        Co2[245]<=(1&0|(1|0)&Co2[244]);

        Sum2[246]<=1^0^Co2[245];
        Co2[246]<=(1&0|(1|0)&Co2[245]);

        Sum2[247]<=1^0^Co2[246];
        Co2[247]<=(1&0|(1|0)&Co2[246]);

        Sum2[248]<=1^0^Co2[247];
        Co2[248]<=(1&0|(1|0)&Co2[247]);

        Sum2[249]<=1^0^Co2[248];
        Co2[249]<=(1&0|(1|0)&Co2[248]);

        Sum2[250]<=1^0^Co2[249];
        Co2[250]<=(1&0|(1|0)&Co2[249]);

        Sum2[251]<=1^0^Co2[250];
        Co2[251]<=(1&0|(1|0)&Co2[250]);

        Sum2[252]<=1^0^Co2[251];
        Co2[252]<=(1&0|(1|0)&Co2[251]);

        Sum2[253]<=1^0^Co2[252];
        Co2[253]<=(1&0|(1|0)&Co2[252]);

        Sum2[254]<=1^0^Co2[253];
        Co2[254]<=(1&0|(1|0)&Co2[253]);

        Sum2[255]<=1^0^Co2[254];
        Co2[255]<=(1&0|(1|0)&Co2[254]);

        Sum2[256]<=1^0^Co2[255];
        Co2[256]<=(1&0|(1|0)&Co2[255]);

        Sum2[257]<=1^0^Co2[256];
        Co2[257]<=(1&0|(1|0)&Co2[256]);

        Sum2[258]<=1^0^Co2[257];
        Co2[258]<=(1&0|(1|0)&Co2[257]);

        Sum2[259]<=1^0^Co2[258];
        Co2[259]<=(1&0|(1|0)&Co2[258]);

        Sum2[260]<=1^0^Co2[259];
        Co2[260]<=(1&0|(1|0)&Co2[259]);

        Sum2[261]<=1^0^Co2[260];
        Co2[261]<=(1&0|(1|0)&Co2[260]);

        Sum2[262]<=1^0^Co2[261];
        Co2[262]<=(1&0|(1|0)&Co2[261]);

        Sum2[263]<=1^0^Co2[262];
        Co2[263]<=(1&0|(1|0)&Co2[262]);

        Sum2[264]<=1^0^Co2[263];
        Co2[264]<=(1&0|(1|0)&Co2[263]);

        Sum2[265]<=1^0^Co2[264];
        Co2[265]<=(1&0|(1|0)&Co2[264]);

        Sum2[266]<=1^0^Co2[265];
        Co2[266]<=(1&0|(1|0)&Co2[265]);

        Sum2[267]<=1^0^Co2[266];
        Co2[267]<=(1&0|(1|0)&Co2[266]);

        Sum2[268]<=1^0^Co2[267];
        Co2[268]<=(1&0|(1|0)&Co2[267]);

        Sum2[269]<=1^0^Co2[268];
        Co2[269]<=(1&0|(1|0)&Co2[268]);

        Sum2[270]<=1^0^Co2[269];
        Co2[270]<=(1&0|(1|0)&Co2[269]);

        Sum2[271]<=1^0^Co2[270];
        Co2[271]<=(1&0|(1|0)&Co2[270]);

        Sum2[272]<=1^0^Co2[271];
        Co2[272]<=(1&0|(1|0)&Co2[271]);

        Sum2[273]<=1^0^Co2[272];
        Co2[273]<=(1&0|(1|0)&Co2[272]);

        Sum2[274]<=1^0^Co2[273];
        Co2[274]<=(1&0|(1|0)&Co2[273]);

        Sum2[275]<=1^0^Co2[274];
        Co2[275]<=(1&0|(1|0)&Co2[274]);

        Sum2[276]<=1^0^Co2[275];
        Co2[276]<=(1&0|(1|0)&Co2[275]);

        Sum2[277]<=1^0^Co2[276];
        Co2[277]<=(1&0|(1|0)&Co2[276]);

        Sum2[278]<=1^0^Co2[277];
        Co2[278]<=(1&0|(1|0)&Co2[277]);

        Sum2[279]<=1^0^Co2[278];
        Co2[279]<=(1&0|(1|0)&Co2[278]);

        Sum2[280]<=1^0^Co2[279];
        Co2[280]<=(1&0|(1|0)&Co2[279]);

        Sum2[281]<=1^0^Co2[280];
        Co2[281]<=(1&0|(1|0)&Co2[280]);

        Sum2[282]<=1^0^Co2[281];
        Co2[282]<=(1&0|(1|0)&Co2[281]);

        Sum2[283]<=1^0^Co2[282];
        Co2[283]<=(1&0|(1|0)&Co2[282]);

        Sum2[284]<=1^0^Co2[283];
        Co2[284]<=(1&0|(1|0)&Co2[283]);

        Sum2[285]<=1^0^Co2[284];
        Co2[285]<=(1&0|(1|0)&Co2[284]);

        Sum2[286]<=1^0^Co2[285];
        Co2[286]<=(1&0|(1|0)&Co2[285]);

        Sum2[287]<=1^0^Co2[286];
        Co2[287]<=(1&0|(1|0)&Co2[286]);

        Sum2[288]<=1^0^Co2[287];
        Co2[288]<=(1&0|(1|0)&Co2[287]);

        Sum2[289]<=1^0^Co2[288];
        Co2[289]<=(1&0|(1|0)&Co2[288]);

        Sum2[290]<=1^0^Co2[289];
        Co2[290]<=(1&0|(1|0)&Co2[289]);

        Sum2[291]<=1^0^Co2[290];
        Co2[291]<=(1&0|(1|0)&Co2[290]);

        Sum2[292]<=1^0^Co2[291];
        Co2[292]<=(1&0|(1|0)&Co2[291]);

        Sum2[293]<=1^0^Co2[292];
        Co2[293]<=(1&0|(1|0)&Co2[292]);

        Sum2[294]<=1^0^Co2[293];
        Co2[294]<=(1&0|(1|0)&Co2[293]);

        Sum2[295]<=1^0^Co2[294];
        Co2[295]<=(1&0|(1|0)&Co2[294]);

        Sum2[296]<=1^0^Co2[295];
        Co2[296]<=(1&0|(1|0)&Co2[295]);

        Sum2[297]<=1^0^Co2[296];
        Co2[297]<=(1&0|(1|0)&Co2[296]);

        Sum2[298]<=1^0^Co2[297];
        Co2[298]<=(1&0|(1|0)&Co2[297]);

        Sum2[299]<=1^0^Co2[298];
        Co2[299]<=(1&0|(1|0)&Co2[298]);

        Sum2[300]<=1^0^Co2[299];
        Co2[300]<=(1&0|(1|0)&Co2[299]);

        Sum2[301]<=1^0^Co2[300];
        Co2[301]<=(1&0|(1|0)&Co2[300]);

        Sum2[302]<=1^0^Co2[301];
        Co2[302]<=(1&0|(1|0)&Co2[301]);

        Sum2[303]<=1^0^Co2[302];
        Co2[303]<=(1&0|(1|0)&Co2[302]);

        Sum2[304]<=1^0^Co2[303];
        Co2[304]<=(1&0|(1|0)&Co2[303]);

        Sum2[305]<=1^0^Co2[304];
        Co2[305]<=(1&0|(1|0)&Co2[304]);

        Sum2[306]<=1^0^Co2[305];
        Co2[306]<=(1&0|(1|0)&Co2[305]);

        Sum2[307]<=1^0^Co2[306];
        Co2[307]<=(1&0|(1|0)&Co2[306]);

        Sum2[308]<=1^0^Co2[307];
        Co2[308]<=(1&0|(1|0)&Co2[307]);

        Sum2[309]<=1^0^Co2[308];
        Co2[309]<=(1&0|(1|0)&Co2[308]);

        Sum2[310]<=1^0^Co2[309];
        Co2[310]<=(1&0|(1|0)&Co2[309]);

        Sum2[311]<=1^0^Co2[310];
        Co2[311]<=(1&0|(1|0)&Co2[310]);

        Sum2[312]<=1^0^Co2[311];
        Co2[312]<=(1&0|(1|0)&Co2[311]);

        Sum2[313]<=1^0^Co2[312];
        Co2[313]<=(1&0|(1|0)&Co2[312]);

        Sum2[314]<=1^0^Co2[313];
        Co2[314]<=(1&0|(1|0)&Co2[313]);

        Sum2[315]<=1^0^Co2[314];
        Co2[315]<=(1&0|(1|0)&Co2[314]);

        Sum2[316]<=1^0^Co2[315];
        Co2[316]<=(1&0|(1|0)&Co2[315]);

        Sum2[317]<=1^0^Co2[316];
        Co2[317]<=(1&0|(1|0)&Co2[316]);

        Sum2[318]<=1^0^Co2[317];
        Co2[318]<=(1&0|(1|0)&Co2[317]);

        Sum2[319]<=1^0^Co2[318];
        Co2[319]<=(1&0|(1|0)&Co2[318]);

        Sum2[320]<=1^0^Co2[319];
        Co2[320]<=(1&0|(1|0)&Co2[319]);

        Sum2[321]<=1^0^Co2[320];
        Co2[321]<=(1&0|(1|0)&Co2[320]);

        Sum2[322]<=1^0^Co2[321];
        Co2[322]<=(1&0|(1|0)&Co2[321]);

        Sum2[323]<=1^0^Co2[322];
        Co2[323]<=(1&0|(1|0)&Co2[322]);

        Sum2[324]<=1^0^Co2[323];
        Co2[324]<=(1&0|(1|0)&Co2[323]);

        Sum2[325]<=1^0^Co2[324];
        Co2[325]<=(1&0|(1|0)&Co2[324]);

        Sum2[326]<=1^0^Co2[325];
        Co2[326]<=(1&0|(1|0)&Co2[325]);

        Sum2[327]<=1^0^Co2[326];
        Co2[327]<=(1&0|(1|0)&Co2[326]);

        Sum2[328]<=1^0^Co2[327];
        Co2[328]<=(1&0|(1|0)&Co2[327]);

        Sum2[329]<=1^0^Co2[328];
        Co2[329]<=(1&0|(1|0)&Co2[328]);

        Sum2[330]<=1^0^Co2[329];
        Co2[330]<=(1&0|(1|0)&Co2[329]);

        Sum2[331]<=1^0^Co2[330];
        Co2[331]<=(1&0|(1|0)&Co2[330]);

        Sum2[332]<=1^0^Co2[331];
        Co2[332]<=(1&0|(1|0)&Co2[331]);

        Sum2[333]<=1^0^Co2[332];
        Co2[333]<=(1&0|(1|0)&Co2[332]);

        Sum2[334]<=1^0^Co2[333];
        Co2[334]<=(1&0|(1|0)&Co2[333]);

        Sum2[335]<=1^0^Co2[334];
        Co2[335]<=(1&0|(1|0)&Co2[334]);

        Sum2[336]<=1^0^Co2[335];
        Co2[336]<=(1&0|(1|0)&Co2[335]);

        Sum2[337]<=1^0^Co2[336];
        Co2[337]<=(1&0|(1|0)&Co2[336]);

        Sum2[338]<=1^0^Co2[337];
        Co2[338]<=(1&0|(1|0)&Co2[337]);

        Sum2[339]<=1^0^Co2[338];
        Co2[339]<=(1&0|(1|0)&Co2[338]);

        Sum2[340]<=1^0^Co2[339];
        Co2[340]<=(1&0|(1|0)&Co2[339]);

        Sum2[341]<=1^0^Co2[340];
        Co2[341]<=(1&0|(1|0)&Co2[340]);

        Sum2[342]<=1^0^Co2[341];
        Co2[342]<=(1&0|(1|0)&Co2[341]);

        Sum2[343]<=1^0^Co2[342];
        Co2[343]<=(1&0|(1|0)&Co2[342]);

        Sum2[344]<=1^0^Co2[343];
        Co2[344]<=(1&0|(1|0)&Co2[343]);

        Sum2[345]<=1^0^Co2[344];
        Co2[345]<=(1&0|(1|0)&Co2[344]);

        Sum2[346]<=1^0^Co2[345];
        Co2[346]<=(1&0|(1|0)&Co2[345]);

        Sum2[347]<=1^0^Co2[346];
        Co2[347]<=(1&0|(1|0)&Co2[346]);

        Sum2[348]<=1^0^Co2[347];
        Co2[348]<=(1&0|(1|0)&Co2[347]);

        Sum2[349]<=1^0^Co2[348];
        Co2[349]<=(1&0|(1|0)&Co2[348]);

        Sum2[350]<=1^0^Co2[349];
        Co2[350]<=(1&0|(1|0)&Co2[349]);

        Sum2[351]<=1^0^Co2[350];
        Co2[351]<=(1&0|(1|0)&Co2[350]);

        Sum2[352]<=1^0^Co2[351];
        Co2[352]<=(1&0|(1|0)&Co2[351]);

        Sum2[353]<=1^0^Co2[352];
        Co2[353]<=(1&0|(1|0)&Co2[352]);

        Sum2[354]<=1^0^Co2[353];
        Co2[354]<=(1&0|(1|0)&Co2[353]);

        Sum2[355]<=1^0^Co2[354];
        Co2[355]<=(1&0|(1|0)&Co2[354]);

        Sum2[356]<=1^0^Co2[355];
        Co2[356]<=(1&0|(1|0)&Co2[355]);

        Sum2[357]<=1^0^Co2[356];
        Co2[357]<=(1&0|(1|0)&Co2[356]);

        Sum2[358]<=1^0^Co2[357];
        Co2[358]<=(1&0|(1|0)&Co2[357]);

        Sum2[359]<=1^0^Co2[358];
        Co2[359]<=(1&0|(1|0)&Co2[358]);

        Sum2[360]<=1^0^Co2[359];
        Co2[360]<=(1&0|(1|0)&Co2[359]);

        Sum2[361]<=1^0^Co2[360];
        Co2[361]<=(1&0|(1|0)&Co2[360]);

        Sum2[362]<=1^0^Co2[361];
        Co2[362]<=(1&0|(1|0)&Co2[361]);

        Sum2[363]<=1^0^Co2[362];
        Co2[363]<=(1&0|(1|0)&Co2[362]);

        Sum2[364]<=1^0^Co2[363];
        Co2[364]<=(1&0|(1|0)&Co2[363]);

        Sum2[365]<=1^0^Co2[364];
        Co2[365]<=(1&0|(1|0)&Co2[364]);

        Sum2[366]<=1^0^Co2[365];
        Co2[366]<=(1&0|(1|0)&Co2[365]);

        Sum2[367]<=1^0^Co2[366];
        Co2[367]<=(1&0|(1|0)&Co2[366]);

        Sum2[368]<=1^0^Co2[367];
        Co2[368]<=(1&0|(1|0)&Co2[367]);

        Sum2[369]<=1^0^Co2[368];
        Co2[369]<=(1&0|(1|0)&Co2[368]);

        Sum2[370]<=1^0^Co2[369];
        Co2[370]<=(1&0|(1|0)&Co2[369]);

        Sum2[371]<=1^0^Co2[370];
        Co2[371]<=(1&0|(1|0)&Co2[370]);

        Sum2[372]<=1^0^Co2[371];
        Co2[372]<=(1&0|(1|0)&Co2[371]);

        Sum2[373]<=1^0^Co2[372];
        Co2[373]<=(1&0|(1|0)&Co2[372]);

        Sum2[374]<=1^0^Co2[373];
        Co2[374]<=(1&0|(1|0)&Co2[373]);

        Sum2[375]<=1^0^Co2[374];
        Co2[375]<=(1&0|(1|0)&Co2[374]);

        Sum2[376]<=1^0^Co2[375];
        Co2[376]<=(1&0|(1|0)&Co2[375]);

        Sum2[377]<=1^0^Co2[376];
        Co2[377]<=(1&0|(1|0)&Co2[376]);

        Sum2[378]<=1^0^Co2[377];
        Co2[378]<=(1&0|(1|0)&Co2[377]);

        Sum2[379]<=1^0^Co2[378];
        Co2[379]<=(1&0|(1|0)&Co2[378]);

        Sum2[380]<=1^0^Co2[379];
        Co2[380]<=(1&0|(1|0)&Co2[379]);

        Sum2[381]<=1^0^Co2[380];
        Co2[381]<=(1&0|(1|0)&Co2[380]);

        Sum2[382]<=1^0^Co2[381];
        Co2[382]<=(1&0|(1|0)&Co2[381]);

        Sum2[383]<=1^0^Co2[382];
        Co2[383]<=(1&0|(1|0)&Co2[382]);

        Sum2[384]<=1^0^Co2[383];
        Co2[384]<=(1&0|(1|0)&Co2[383]);

        Sum2[385]<=1^0^Co2[384];
        Co2[385]<=(1&0|(1|0)&Co2[384]);

        Sum2[386]<=1^0^Co2[385];
        Co2[386]<=(1&0|(1|0)&Co2[385]);

        Sum2[387]<=1^0^Co2[386];
        Co2[387]<=(1&0|(1|0)&Co2[386]);

        Sum2[388]<=1^0^Co2[387];
        Co2[388]<=(1&0|(1|0)&Co2[387]);

        Sum2[389]<=1^0^Co2[388];
        Co2[389]<=(1&0|(1|0)&Co2[388]);

        Sum2[390]<=1^0^Co2[389];
        Co2[390]<=(1&0|(1|0)&Co2[389]);

        Sum2[391]<=1^0^Co2[390];
        Co2[391]<=(1&0|(1|0)&Co2[390]);

        Sum2[392]<=1^0^Co2[391];
        Co2[392]<=(1&0|(1|0)&Co2[391]);

        Sum2[393]<=1^0^Co2[392];
        Co2[393]<=(1&0|(1|0)&Co2[392]);

        Sum2[394]<=1^0^Co2[393];
        Co2[394]<=(1&0|(1|0)&Co2[393]);

        Sum2[395]<=1^0^Co2[394];
        Co2[395]<=(1&0|(1|0)&Co2[394]);

        Sum2[396]<=1^0^Co2[395];
        Co2[396]<=(1&0|(1|0)&Co2[395]);

        Sum2[397]<=1^0^Co2[396];
        Co2[397]<=(1&0|(1|0)&Co2[396]);

        Sum2[398]<=1^0^Co2[397];
        Co2[398]<=(1&0|(1|0)&Co2[397]);

        Sum2[399]<=1^0^Co2[398];
        Co2[399]<=(1&0|(1|0)&Co2[398]);

        Sum2[400]<=1^0^Co2[399];
        Co2[400]<=(1&0|(1|0)&Co2[399]);

        Sum2[401]<=1^0^Co2[400];
        Co2[401]<=(1&0|(1|0)&Co2[400]);

        Sum2[402]<=1^0^Co2[401];
        Co2[402]<=(1&0|(1|0)&Co2[401]);

        Sum2[403]<=1^0^Co2[402];
        Co2[403]<=(1&0|(1|0)&Co2[402]);

        Sum2[404]<=1^0^Co2[403];
        Co2[404]<=(1&0|(1|0)&Co2[403]);

        Sum2[405]<=1^0^Co2[404];
        Co2[405]<=(1&0|(1|0)&Co2[404]);

        Sum2[406]<=1^0^Co2[405];
        Co2[406]<=(1&0|(1|0)&Co2[405]);

        Sum2[407]<=1^0^Co2[406];
        Co2[407]<=(1&0|(1|0)&Co2[406]);

        Sum2[408]<=1^0^Co2[407];
        Co2[408]<=(1&0|(1|0)&Co2[407]);

        Sum2[409]<=1^0^Co2[408];
        Co2[409]<=(1&0|(1|0)&Co2[408]);

        Sum2[410]<=1^0^Co2[409];
        Co2[410]<=(1&0|(1|0)&Co2[409]);

        Sum2[411]<=1^0^Co2[410];
        Co2[411]<=(1&0|(1|0)&Co2[410]);

        Sum2[412]<=1^0^Co2[411];
        Co2[412]<=(1&0|(1|0)&Co2[411]);

        Sum2[413]<=1^0^Co2[412];
        Co2[413]<=(1&0|(1|0)&Co2[412]);

        Sum2[414]<=1^0^Co2[413];
        Co2[414]<=(1&0|(1|0)&Co2[413]);

        Sum2[415]<=1^0^Co2[414];
        Co2[415]<=(1&0|(1|0)&Co2[414]);

        Sum2[416]<=1^0^Co2[415];
        Co2[416]<=(1&0|(1|0)&Co2[415]);

        Sum2[417]<=1^0^Co2[416];
        Co2[417]<=(1&0|(1|0)&Co2[416]);

        Sum2[418]<=1^0^Co2[417];
        Co2[418]<=(1&0|(1|0)&Co2[417]);

        Sum2[419]<=1^0^Co2[418];
        Co2[419]<=(1&0|(1|0)&Co2[418]);

        Sum2[420]<=1^0^Co2[419];
        Co2[420]<=(1&0|(1|0)&Co2[419]);

        Sum2[421]<=1^0^Co2[420];
        Co2[421]<=(1&0|(1|0)&Co2[420]);

        Sum2[422]<=1^0^Co2[421];
        Co2[422]<=(1&0|(1|0)&Co2[421]);

        Sum2[423]<=1^0^Co2[422];
        Co2[423]<=(1&0|(1|0)&Co2[422]);

        Sum2[424]<=1^0^Co2[423];
        Co2[424]<=(1&0|(1|0)&Co2[423]);

        Sum2[425]<=1^0^Co2[424];
        Co2[425]<=(1&0|(1|0)&Co2[424]);

        Sum2[426]<=1^0^Co2[425];
        Co2[426]<=(1&0|(1|0)&Co2[425]);

        Sum2[427]<=1^0^Co2[426];
        Co2[427]<=(1&0|(1|0)&Co2[426]);

        Sum2[428]<=1^0^Co2[427];
        Co2[428]<=(1&0|(1|0)&Co2[427]);

        Sum2[429]<=1^0^Co2[428];
        Co2[429]<=(1&0|(1|0)&Co2[428]);

        Sum2[430]<=1^0^Co2[429];
        Co2[430]<=(1&0|(1|0)&Co2[429]);

        Sum2[431]<=1^0^Co2[430];
        Co2[431]<=(1&0|(1|0)&Co2[430]);

        Sum2[432]<=1^0^Co2[431];
        Co2[432]<=(1&0|(1|0)&Co2[431]);

        Sum2[433]<=1^0^Co2[432];
        Co2[433]<=(1&0|(1|0)&Co2[432]);

        Sum2[434]<=1^0^Co2[433];
        Co2[434]<=(1&0|(1|0)&Co2[433]);

        Sum2[435]<=1^0^Co2[434];
        Co2[435]<=(1&0|(1|0)&Co2[434]);

        Sum2[436]<=1^0^Co2[435];
        Co2[436]<=(1&0|(1|0)&Co2[435]);

        Sum2[437]<=1^0^Co2[436];
        Co2[437]<=(1&0|(1|0)&Co2[436]);

        Sum2[438]<=1^0^Co2[437];
        Co2[438]<=(1&0|(1|0)&Co2[437]);

        Sum2[439]<=1^0^Co2[438];
        Co2[439]<=(1&0|(1|0)&Co2[438]);

        Sum2[440]<=1^0^Co2[439];
        Co2[440]<=(1&0|(1|0)&Co2[439]);

        Sum2[441]<=1^0^Co2[440];
        Co2[441]<=(1&0|(1|0)&Co2[440]);

        Sum2[442]<=1^0^Co2[441];
        Co2[442]<=(1&0|(1|0)&Co2[441]);

        Sum2[443]<=1^0^Co2[442];
        Co2[443]<=(1&0|(1|0)&Co2[442]);

        Sum2[444]<=1^0^Co2[443];
        Co2[444]<=(1&0|(1|0)&Co2[443]);

        Sum2[445]<=1^0^Co2[444];
        Co2[445]<=(1&0|(1|0)&Co2[444]);

        Sum2[446]<=1^0^Co2[445];
        Co2[446]<=(1&0|(1|0)&Co2[445]);

        Sum2[447]<=1^0^Co2[446];
        Co2[447]<=(1&0|(1|0)&Co2[446]);

        Sum2[448]<=1^0^Co2[447];
        Co2[448]<=(1&0|(1|0)&Co2[447]);

        Sum2[449]<=1^0^Co2[448];
        Co2[449]<=(1&0|(1|0)&Co2[448]);

        Sum2[450]<=1^0^Co2[449];
        Co2[450]<=(1&0|(1|0)&Co2[449]);

        Sum2[451]<=1^0^Co2[450];
        Co2[451]<=(1&0|(1|0)&Co2[450]);

        Sum2[452]<=1^0^Co2[451];
        Co2[452]<=(1&0|(1|0)&Co2[451]);

        Sum2[453]<=1^0^Co2[452];
        Co2[453]<=(1&0|(1|0)&Co2[452]);

        Sum2[454]<=1^0^Co2[453];
        Co2[454]<=(1&0|(1|0)&Co2[453]);

        Sum2[455]<=1^0^Co2[454];
        Co2[455]<=(1&0|(1|0)&Co2[454]);

        Sum2[456]<=1^0^Co2[455];
        Co2[456]<=(1&0|(1|0)&Co2[455]);

        Sum2[457]<=1^0^Co2[456];
        Co2[457]<=(1&0|(1|0)&Co2[456]);

        Sum2[458]<=1^0^Co2[457];
        Co2[458]<=(1&0|(1|0)&Co2[457]);

        Sum2[459]<=1^0^Co2[458];
        Co2[459]<=(1&0|(1|0)&Co2[458]);

        Sum2[460]<=1^0^Co2[459];
        Co2[460]<=(1&0|(1|0)&Co2[459]);

        Sum2[461]<=1^0^Co2[460];
        Co2[461]<=(1&0|(1|0)&Co2[460]);

        Sum2[462]<=1^0^Co2[461];
        Co2[462]<=(1&0|(1|0)&Co2[461]);

        Sum2[463]<=1^0^Co2[462];
        Co2[463]<=(1&0|(1|0)&Co2[462]);

        Sum2[464]<=1^0^Co2[463];
        Co2[464]<=(1&0|(1|0)&Co2[463]);

        Sum2[465]<=1^0^Co2[464];
        Co2[465]<=(1&0|(1|0)&Co2[464]);

        Sum2[466]<=1^0^Co2[465];
        Co2[466]<=(1&0|(1|0)&Co2[465]);

        Sum2[467]<=1^0^Co2[466];
        Co2[467]<=(1&0|(1|0)&Co2[466]);

        Sum2[468]<=1^0^Co2[467];
        Co2[468]<=(1&0|(1|0)&Co2[467]);

        Sum2[469]<=1^0^Co2[468];
        Co2[469]<=(1&0|(1|0)&Co2[468]);

        Sum2[470]<=1^0^Co2[469];
        Co2[470]<=(1&0|(1|0)&Co2[469]);

        Sum2[471]<=1^0^Co2[470];
        Co2[471]<=(1&0|(1|0)&Co2[470]);

        Sum2[472]<=1^0^Co2[471];
        Co2[472]<=(1&0|(1|0)&Co2[471]);

        Sum2[473]<=1^0^Co2[472];
        Co2[473]<=(1&0|(1|0)&Co2[472]);

        Sum2[474]<=1^0^Co2[473];
        Co2[474]<=(1&0|(1|0)&Co2[473]);

        Sum2[475]<=1^0^Co2[474];
        Co2[475]<=(1&0|(1|0)&Co2[474]);

        Sum2[476]<=1^0^Co2[475];
        Co2[476]<=(1&0|(1|0)&Co2[475]);

        Sum2[477]<=1^0^Co2[476];
        Co2[477]<=(1&0|(1|0)&Co2[476]);

        Sum2[478]<=1^0^Co2[477];
        Co2[478]<=(1&0|(1|0)&Co2[477]);

        Sum2[479]<=1^0^Co2[478];
        Co2[479]<=(1&0|(1|0)&Co2[478]);

        Sum2[480]<=1^0^Co2[479];
        Co2[480]<=(1&0|(1|0)&Co2[479]);

        Sum2[481]<=1^0^Co2[480];
        Co2[481]<=(1&0|(1|0)&Co2[480]);

        Sum2[482]<=1^0^Co2[481];
        Co2[482]<=(1&0|(1|0)&Co2[481]);

        Sum2[483]<=1^0^Co2[482];
        Co2[483]<=(1&0|(1|0)&Co2[482]);

        Sum2[484]<=1^0^Co2[483];
        Co2[484]<=(1&0|(1|0)&Co2[483]);

        Sum2[485]<=1^0^Co2[484];
        Co2[485]<=(1&0|(1|0)&Co2[484]);

        Sum2[486]<=1^0^Co2[485];
        Co2[486]<=(1&0|(1|0)&Co2[485]);

        Sum2[487]<=1^0^Co2[486];
        Co2[487]<=(1&0|(1|0)&Co2[486]);

        Sum2[488]<=1^0^Co2[487];
        Co2[488]<=(1&0|(1|0)&Co2[487]);

        Sum2[489]<=1^0^Co2[488];
        Co2[489]<=(1&0|(1|0)&Co2[488]);

        Sum2[490]<=1^0^Co2[489];
        Co2[490]<=(1&0|(1|0)&Co2[489]);

        Sum2[491]<=1^0^Co2[490];
        Co2[491]<=(1&0|(1|0)&Co2[490]);

        Sum2[492]<=1^0^Co2[491];
        Co2[492]<=(1&0|(1|0)&Co2[491]);

        Sum2[493]<=1^0^Co2[492];
        Co2[493]<=(1&0|(1|0)&Co2[492]);

        Sum2[494]<=1^0^Co2[493];
        Co2[494]<=(1&0|(1|0)&Co2[493]);

        Sum2[495]<=1^0^Co2[494];
        Co2[495]<=(1&0|(1|0)&Co2[494]);

        Sum2[496]<=1^0^Co2[495];
        Co2[496]<=(1&0|(1|0)&Co2[495]);

        Sum2[497]<=1^0^Co2[496];
        Co2[497]<=(1&0|(1|0)&Co2[496]);

        Sum2[498]<=1^0^Co2[497];
        Co2[498]<=(1&0|(1|0)&Co2[497]);

        Sum2[499]<=1^0^Co2[498];
        Co2[499]<=(1&0|(1|0)&Co2[498]);

        Sum2[500]<=1^0^Co2[499];
        Co2[500]<=(1&0|(1|0)&Co2[499]);

        Sum2[501]<=1^0^Co2[500];
        Co2[501]<=(1&0|(1|0)&Co2[500]);

        Sum2[502]<=1^0^Co2[501];
        Co2[502]<=(1&0|(1|0)&Co2[501]);

        Sum2[503]<=1^0^Co2[502];
        Co2[503]<=(1&0|(1|0)&Co2[502]);

        Sum2[504]<=1^0^Co2[503];
        Co2[504]<=(1&0|(1|0)&Co2[503]);

        Sum2[505]<=1^0^Co2[504];
        Co2[505]<=(1&0|(1|0)&Co2[504]);

        Sum2[506]<=1^0^Co2[505];
        Co2[506]<=(1&0|(1|0)&Co2[505]);

        Sum2[507]<=1^0^Co2[506];
        Co2[507]<=(1&0|(1|0)&Co2[506]);

        Sum2[508]<=1^0^Co2[507];
        Co2[508]<=(1&0|(1|0)&Co2[507]);

        Sum2[509]<=1^0^Co2[508];
        Co2[509]<=(1&0|(1|0)&Co2[508]);

        Sum2[510]<=1^0^Co2[509];
        Co2[510]<=(1&0|(1|0)&Co2[509]);

        Sum2[511]<=1^0^Co2[510];
        Co2[511]<=(1&0|(1|0)&Co2[510]);

        Sum2[512]<=1^0^Co2[511];
        Co2[512]<=(1&0|(1|0)&Co2[511]);

        Sum2[513]<=1^0^Co2[512];
        Co2[513]<=(1&0|(1|0)&Co2[512]);

        Sum2[514]<=1^0^Co2[513];
        Co2[514]<=(1&0|(1|0)&Co2[513]);

        Sum2[515]<=1^0^Co2[514];
        Co2[515]<=(1&0|(1|0)&Co2[514]);

        Sum2[516]<=1^0^Co2[515];
        Co2[516]<=(1&0|(1|0)&Co2[515]);

        Sum2[517]<=1^0^Co2[516];
        Co2[517]<=(1&0|(1|0)&Co2[516]);

        Sum2[518]<=1^0^Co2[517];
        Co2[518]<=(1&0|(1|0)&Co2[517]);

        Sum2[519]<=1^0^Co2[518];
        Co2[519]<=(1&0|(1|0)&Co2[518]);

        Sum2[520]<=1^0^Co2[519];
        Co2[520]<=(1&0|(1|0)&Co2[519]);

        Sum2[521]<=1^0^Co2[520];
        Co2[521]<=(1&0|(1|0)&Co2[520]);

        Sum2[522]<=1^0^Co2[521];
        Co2[522]<=(1&0|(1|0)&Co2[521]);

        Sum2[523]<=1^0^Co2[522];
        Co2[523]<=(1&0|(1|0)&Co2[522]);

        Sum2[524]<=1^0^Co2[523];
        Co2[524]<=(1&0|(1|0)&Co2[523]);

        Sum2[525]<=1^0^Co2[524];
        Co2[525]<=(1&0|(1|0)&Co2[524]);

        Sum2[526]<=1^0^Co2[525];
        Co2[526]<=(1&0|(1|0)&Co2[525]);

        Sum2[527]<=1^0^Co2[526];
        Co2[527]<=(1&0|(1|0)&Co2[526]);

        Sum2[528]<=1^0^Co2[527];
        Co2[528]<=(1&0|(1|0)&Co2[527]);

        Sum2[529]<=1^0^Co2[528];
        Co2[529]<=(1&0|(1|0)&Co2[528]);

        Sum2[530]<=1^0^Co2[529];
        Co2[530]<=(1&0|(1|0)&Co2[529]);

        Sum2[531]<=1^0^Co2[530];
        Co2[531]<=(1&0|(1|0)&Co2[530]);

        Sum2[532]<=1^0^Co2[531];
        Co2[532]<=(1&0|(1|0)&Co2[531]);

        Sum2[533]<=1^0^Co2[532];
        Co2[533]<=(1&0|(1|0)&Co2[532]);

        Sum2[534]<=1^0^Co2[533];
        Co2[534]<=(1&0|(1|0)&Co2[533]);

        Sum2[535]<=1^0^Co2[534];
        Co2[535]<=(1&0|(1|0)&Co2[534]);

        Sum2[536]<=1^0^Co2[535];
        Co2[536]<=(1&0|(1|0)&Co2[535]);

        Sum2[537]<=1^0^Co2[536];
        Co2[537]<=(1&0|(1|0)&Co2[536]);

        Sum2[538]<=1^0^Co2[537];
        Co2[538]<=(1&0|(1|0)&Co2[537]);

        Sum2[539]<=1^0^Co2[538];
        Co2[539]<=(1&0|(1|0)&Co2[538]);

        Sum2[540]<=1^0^Co2[539];
        Co2[540]<=(1&0|(1|0)&Co2[539]);

        Sum2[541]<=1^0^Co2[540];
        Co2[541]<=(1&0|(1|0)&Co2[540]);

        Sum2[542]<=1^0^Co2[541];
        Co2[542]<=(1&0|(1|0)&Co2[541]);

        Sum2[543]<=1^0^Co2[542];
        Co2[543]<=(1&0|(1|0)&Co2[542]);

        Sum2[544]<=1^0^Co2[543];
        Co2[544]<=(1&0|(1|0)&Co2[543]);

        Sum2[545]<=1^0^Co2[544];
        Co2[545]<=(1&0|(1|0)&Co2[544]);

        Sum2[546]<=1^0^Co2[545];
        Co2[546]<=(1&0|(1|0)&Co2[545]);

        Sum2[547]<=1^0^Co2[546];
        Co2[547]<=(1&0|(1|0)&Co2[546]);

        Sum2[548]<=1^0^Co2[547];
        Co2[548]<=(1&0|(1|0)&Co2[547]);

        Sum2[549]<=1^0^Co2[548];
        Co2[549]<=(1&0|(1|0)&Co2[548]);

        Sum2[550]<=1^0^Co2[549];
        Co2[550]<=(1&0|(1|0)&Co2[549]);

        Sum2[551]<=1^0^Co2[550];
        Co2[551]<=(1&0|(1|0)&Co2[550]);

        Sum2[552]<=1^0^Co2[551];
        Co2[552]<=(1&0|(1|0)&Co2[551]);

        Sum2[553]<=1^0^Co2[552];
        Co2[553]<=(1&0|(1|0)&Co2[552]);

        Sum2[554]<=1^0^Co2[553];
        Co2[554]<=(1&0|(1|0)&Co2[553]);

        Sum2[555]<=1^0^Co2[554];
        Co2[555]<=(1&0|(1|0)&Co2[554]);

        Sum2[556]<=1^0^Co2[555];
        Co2[556]<=(1&0|(1|0)&Co2[555]);

        Sum2[557]<=1^0^Co2[556];
        Co2[557]<=(1&0|(1|0)&Co2[556]);

        Sum2[558]<=1^0^Co2[557];
        Co2[558]<=(1&0|(1|0)&Co2[557]);

        Sum2[559]<=1^0^Co2[558];
        Co2[559]<=(1&0|(1|0)&Co2[558]);

        Sum2[560]<=1^0^Co2[559];
        Co2[560]<=(1&0|(1|0)&Co2[559]);

        Sum2[561]<=1^0^Co2[560];
        Co2[561]<=(1&0|(1|0)&Co2[560]);

        Sum2[562]<=1^0^Co2[561];
        Co2[562]<=(1&0|(1|0)&Co2[561]);

        Sum2[563]<=1^0^Co2[562];
        Co2[563]<=(1&0|(1|0)&Co2[562]);

        Sum2[564]<=1^0^Co2[563];
        Co2[564]<=(1&0|(1|0)&Co2[563]);

        Sum2[565]<=1^0^Co2[564];
        Co2[565]<=(1&0|(1|0)&Co2[564]);

        Sum2[566]<=1^0^Co2[565];
        Co2[566]<=(1&0|(1|0)&Co2[565]);

        Sum2[567]<=1^0^Co2[566];
        Co2[567]<=(1&0|(1|0)&Co2[566]);

        Sum2[568]<=1^0^Co2[567];
        Co2[568]<=(1&0|(1|0)&Co2[567]);

        Sum2[569]<=1^0^Co2[568];
        Co2[569]<=(1&0|(1|0)&Co2[568]);

        Sum2[570]<=1^0^Co2[569];
        Co2[570]<=(1&0|(1|0)&Co2[569]);

        Sum2[571]<=1^0^Co2[570];
        Co2[571]<=(1&0|(1|0)&Co2[570]);

        Sum2[572]<=1^0^Co2[571];
        Co2[572]<=(1&0|(1|0)&Co2[571]);

        Sum2[573]<=1^0^Co2[572];
        Co2[573]<=(1&0|(1|0)&Co2[572]);

        Sum2[574]<=1^0^Co2[573];
        Co2[574]<=(1&0|(1|0)&Co2[573]);

        Sum2[575]<=1^0^Co2[574];
        Co2[575]<=(1&0|(1|0)&Co2[574]);

        Sum2[576]<=1^0^Co2[575];
        Co2[576]<=(1&0|(1|0)&Co2[575]);

        Sum2[577]<=1^0^Co2[576];
        Co2[577]<=(1&0|(1|0)&Co2[576]);

        Sum2[578]<=1^0^Co2[577];
        Co2[578]<=(1&0|(1|0)&Co2[577]);

        Sum2[579]<=1^0^Co2[578];
        Co2[579]<=(1&0|(1|0)&Co2[578]);

        Sum2[580]<=1^0^Co2[579];
        Co2[580]<=(1&0|(1|0)&Co2[579]);

        Sum2[581]<=1^0^Co2[580];
        Co2[581]<=(1&0|(1|0)&Co2[580]);

        Sum2[582]<=1^0^Co2[581];
        Co2[582]<=(1&0|(1|0)&Co2[581]);

        Sum2[583]<=1^0^Co2[582];
        Co2[583]<=(1&0|(1|0)&Co2[582]);

        Sum2[584]<=1^0^Co2[583];
        Co2[584]<=(1&0|(1|0)&Co2[583]);

        Sum2[585]<=1^0^Co2[584];
        Co2[585]<=(1&0|(1|0)&Co2[584]);

        Sum2[586]<=1^0^Co2[585];
        Co2[586]<=(1&0|(1|0)&Co2[585]);

        Sum2[587]<=1^0^Co2[586];
        Co2[587]<=(1&0|(1|0)&Co2[586]);

        Sum2[588]<=1^0^Co2[587];
        Co2[588]<=(1&0|(1|0)&Co2[587]);

        Sum2[589]<=1^0^Co2[588];
        Co2[589]<=(1&0|(1|0)&Co2[588]);

        Sum2[590]<=1^0^Co2[589];
        Co2[590]<=(1&0|(1|0)&Co2[589]);

        Sum2[591]<=1^0^Co2[590];
        Co2[591]<=(1&0|(1|0)&Co2[590]);

        Sum2[592]<=1^0^Co2[591];
        Co2[592]<=(1&0|(1|0)&Co2[591]);

        Sum2[593]<=1^0^Co2[592];
        Co2[593]<=(1&0|(1|0)&Co2[592]);

        Sum2[594]<=1^0^Co2[593];
        Co2[594]<=(1&0|(1|0)&Co2[593]);

        Sum2[595]<=1^0^Co2[594];
        Co2[595]<=(1&0|(1|0)&Co2[594]);

        Sum2[596]<=1^0^Co2[595];
        Co2[596]<=(1&0|(1|0)&Co2[595]);

        Sum2[597]<=1^0^Co2[596];
        Co2[597]<=(1&0|(1|0)&Co2[596]);

        Sum2[598]<=1^0^Co2[597];
        Co2[598]<=(1&0|(1|0)&Co2[597]);

        Sum2[599]<=1^0^Co2[598];
        Co2[599]<=(1&0|(1|0)&Co2[598]);

        Sum2[600]<=1^0^Co2[599];
        Co2[600]<=(1&0|(1|0)&Co2[599]);

        Sum2[601]<=1^0^Co2[600];
        Co2[601]<=(1&0|(1|0)&Co2[600]);

        Sum2[602]<=1^0^Co2[601];
        Co2[602]<=(1&0|(1|0)&Co2[601]);

        Sum2[603]<=1^0^Co2[602];
        Co2[603]<=(1&0|(1|0)&Co2[602]);

        Sum2[604]<=1^0^Co2[603];
        Co2[604]<=(1&0|(1|0)&Co2[603]);

        Sum2[605]<=1^0^Co2[604];
        Co2[605]<=(1&0|(1|0)&Co2[604]);

        Sum2[606]<=1^0^Co2[605];
        Co2[606]<=(1&0|(1|0)&Co2[605]);

        Sum2[607]<=1^0^Co2[606];
        Co2[607]<=(1&0|(1|0)&Co2[606]);

        Sum2[608]<=1^0^Co2[607];
        Co2[608]<=(1&0|(1|0)&Co2[607]);

        Sum2[609]<=1^0^Co2[608];
        Co2[609]<=(1&0|(1|0)&Co2[608]);

        Sum2[610]<=1^0^Co2[609];
        Co2[610]<=(1&0|(1|0)&Co2[609]);

        Sum2[611]<=1^0^Co2[610];
        Co2[611]<=(1&0|(1|0)&Co2[610]);

        Sum2[612]<=1^0^Co2[611];
        Co2[612]<=(1&0|(1|0)&Co2[611]);

        Sum2[613]<=1^0^Co2[612];
        Co2[613]<=(1&0|(1|0)&Co2[612]);

        Sum2[614]<=1^0^Co2[613];
        Co2[614]<=(1&0|(1|0)&Co2[613]);

        Sum2[615]<=1^0^Co2[614];
        Co2[615]<=(1&0|(1|0)&Co2[614]);

        Sum2[616]<=1^0^Co2[615];
        Co2[616]<=(1&0|(1|0)&Co2[615]);

        Sum2[617]<=1^0^Co2[616];
        Co2[617]<=(1&0|(1|0)&Co2[616]);

        Sum2[618]<=1^0^Co2[617];
        Co2[618]<=(1&0|(1|0)&Co2[617]);

        Sum2[619]<=1^0^Co2[618];
        Co2[619]<=(1&0|(1|0)&Co2[618]);

        Sum2[620]<=1^0^Co2[619];
        Co2[620]<=(1&0|(1|0)&Co2[619]);

        Sum2[621]<=1^0^Co2[620];
        Co2[621]<=(1&0|(1|0)&Co2[620]);

        Sum2[622]<=1^0^Co2[621];
        Co2[622]<=(1&0|(1|0)&Co2[621]);

        Sum2[623]<=1^0^Co2[622];
        Co2[623]<=(1&0|(1|0)&Co2[622]);

        Sum2[624]<=1^0^Co2[623];
        Co2[624]<=(1&0|(1|0)&Co2[623]);

        Sum2[625]<=1^0^Co2[624];
        Co2[625]<=(1&0|(1|0)&Co2[624]);

        Sum2[626]<=1^0^Co2[625];
        Co2[626]<=(1&0|(1|0)&Co2[625]);

        Sum2[627]<=1^0^Co2[626];
        Co2[627]<=(1&0|(1|0)&Co2[626]);

        Sum2[628]<=1^0^Co2[627];
        Co2[628]<=(1&0|(1|0)&Co2[627]);

        Sum2[629]<=1^0^Co2[628];
        Co2[629]<=(1&0|(1|0)&Co2[628]);

        Sum2[630]<=1^0^Co2[629];
        Co2[630]<=(1&0|(1|0)&Co2[629]);

        Sum2[631]<=1^0^Co2[630];
        Co2[631]<=(1&0|(1|0)&Co2[630]);

        Sum2[632]<=1^0^Co2[631];
        Co2[632]<=(1&0|(1|0)&Co2[631]);

        Sum2[633]<=1^0^Co2[632];
        Co2[633]<=(1&0|(1|0)&Co2[632]);

        Sum2[634]<=1^0^Co2[633];
        Co2[634]<=(1&0|(1|0)&Co2[633]);

        Sum2[635]<=1^0^Co2[634];
        Co2[635]<=(1&0|(1|0)&Co2[634]);

        Sum2[636]<=1^0^Co2[635];
        Co2[636]<=(1&0|(1|0)&Co2[635]);

        Sum2[637]<=1^0^Co2[636];
        Co2[637]<=(1&0|(1|0)&Co2[636]);

        Sum2[638]<=1^0^Co2[637];
        Co2[638]<=(1&0|(1|0)&Co2[637]);

        Sum2[639]<=1^0^Co2[638];
        Co2[639]<=(1&0|(1|0)&Co2[638]);

        Sum2[640]<=1^0^Co2[639];
        Co2[640]<=(1&0|(1|0)&Co2[639]);

        Sum2[641]<=1^0^Co2[640];
        Co2[641]<=(1&0|(1|0)&Co2[640]);

        Sum2[642]<=1^0^Co2[641];
        Co2[642]<=(1&0|(1|0)&Co2[641]);

        Sum2[643]<=1^0^Co2[642];
        Co2[643]<=(1&0|(1|0)&Co2[642]);

        Sum2[644]<=1^0^Co2[643];
        Co2[644]<=(1&0|(1|0)&Co2[643]);

        Sum2[645]<=1^0^Co2[644];
        Co2[645]<=(1&0|(1|0)&Co2[644]);

        Sum2[646]<=1^0^Co2[645];
        Co2[646]<=(1&0|(1|0)&Co2[645]);

        Sum2[647]<=1^0^Co2[646];
        Co2[647]<=(1&0|(1|0)&Co2[646]);

        Sum2[648]<=1^0^Co2[647];
        Co2[648]<=(1&0|(1|0)&Co2[647]);

        Sum2[649]<=1^0^Co2[648];
        Co2[649]<=(1&0|(1|0)&Co2[648]);

        Sum2[650]<=1^0^Co2[649];
        Co2[650]<=(1&0|(1|0)&Co2[649]);

        Sum2[651]<=1^0^Co2[650];
        Co2[651]<=(1&0|(1|0)&Co2[650]);

        Sum2[652]<=1^0^Co2[651];
        Co2[652]<=(1&0|(1|0)&Co2[651]);

        Sum2[653]<=1^0^Co2[652];
        Co2[653]<=(1&0|(1|0)&Co2[652]);

        Sum2[654]<=1^0^Co2[653];
        Co2[654]<=(1&0|(1|0)&Co2[653]);

        Sum2[655]<=1^0^Co2[654];
        Co2[655]<=(1&0|(1|0)&Co2[654]);

        Sum2[656]<=1^0^Co2[655];
        Co2[656]<=(1&0|(1|0)&Co2[655]);

        Sum2[657]<=1^0^Co2[656];
        Co2[657]<=(1&0|(1|0)&Co2[656]);

        Sum2[658]<=1^0^Co2[657];
        Co2[658]<=(1&0|(1|0)&Co2[657]);

        Sum2[659]<=1^0^Co2[658];
        Co2[659]<=(1&0|(1|0)&Co2[658]);

        Sum2[660]<=1^0^Co2[659];
        Co2[660]<=(1&0|(1|0)&Co2[659]);

        Sum2[661]<=1^0^Co2[660];
        Co2[661]<=(1&0|(1|0)&Co2[660]);

        Sum2[662]<=1^0^Co2[661];
        Co2[662]<=(1&0|(1|0)&Co2[661]);

        Sum2[663]<=1^0^Co2[662];
        Co2[663]<=(1&0|(1|0)&Co2[662]);

        Sum2[664]<=1^0^Co2[663];
        Co2[664]<=(1&0|(1|0)&Co2[663]);

        Sum2[665]<=1^0^Co2[664];
        Co2[665]<=(1&0|(1|0)&Co2[664]);

        Sum2[666]<=1^0^Co2[665];
        Co2[666]<=(1&0|(1|0)&Co2[665]);

        Sum2[667]<=1^0^Co2[666];
        Co2[667]<=(1&0|(1|0)&Co2[666]);

        Sum2[668]<=1^0^Co2[667];
        Co2[668]<=(1&0|(1|0)&Co2[667]);

        Sum2[669]<=1^0^Co2[668];
        Co2[669]<=(1&0|(1|0)&Co2[668]);

        Sum2[670]<=1^0^Co2[669];
        Co2[670]<=(1&0|(1|0)&Co2[669]);

        Sum2[671]<=1^0^Co2[670];
        Co2[671]<=(1&0|(1|0)&Co2[670]);

        Sum2[672]<=1^0^Co2[671];
        Co2[672]<=(1&0|(1|0)&Co2[671]);

        Sum2[673]<=1^0^Co2[672];
        Co2[673]<=(1&0|(1|0)&Co2[672]);

        Sum2[674]<=1^0^Co2[673];
        Co2[674]<=(1&0|(1|0)&Co2[673]);

        Sum2[675]<=1^0^Co2[674];
        Co2[675]<=(1&0|(1|0)&Co2[674]);

        Sum2[676]<=1^0^Co2[675];
        Co2[676]<=(1&0|(1|0)&Co2[675]);

        Sum2[677]<=1^0^Co2[676];
        Co2[677]<=(1&0|(1|0)&Co2[676]);

        Sum2[678]<=1^0^Co2[677];
        Co2[678]<=(1&0|(1|0)&Co2[677]);

        Sum2[679]<=1^0^Co2[678];
        Co2[679]<=(1&0|(1|0)&Co2[678]);

        Sum2[680]<=1^0^Co2[679];
        Co2[680]<=(1&0|(1|0)&Co2[679]);

        Sum2[681]<=1^0^Co2[680];
        Co2[681]<=(1&0|(1|0)&Co2[680]);

        Sum2[682]<=1^0^Co2[681];
        Co2[682]<=(1&0|(1|0)&Co2[681]);

        Sum2[683]<=1^0^Co2[682];
        Co2[683]<=(1&0|(1|0)&Co2[682]);

        Sum2[684]<=1^0^Co2[683];
        Co2[684]<=(1&0|(1|0)&Co2[683]);

        Sum2[685]<=1^0^Co2[684];
        Co2[685]<=(1&0|(1|0)&Co2[684]);

        Sum2[686]<=1^0^Co2[685];
        Co2[686]<=(1&0|(1|0)&Co2[685]);

        Sum2[687]<=1^0^Co2[686];
        Co2[687]<=(1&0|(1|0)&Co2[686]);

        Sum2[688]<=1^0^Co2[687];
        Co2[688]<=(1&0|(1|0)&Co2[687]);

        Sum2[689]<=1^0^Co2[688];
        Co2[689]<=(1&0|(1|0)&Co2[688]);

        Sum2[690]<=1^0^Co2[689];
        Co2[690]<=(1&0|(1|0)&Co2[689]);

        Sum2[691]<=1^0^Co2[690];
        Co2[691]<=(1&0|(1|0)&Co2[690]);

        Sum2[692]<=1^0^Co2[691];
        Co2[692]<=(1&0|(1|0)&Co2[691]);

        Sum2[693]<=1^0^Co2[692];
        Co2[693]<=(1&0|(1|0)&Co2[692]);

        Sum2[694]<=1^0^Co2[693];
        Co2[694]<=(1&0|(1|0)&Co2[693]);

        Sum2[695]<=1^0^Co2[694];
        Co2[695]<=(1&0|(1|0)&Co2[694]);

        Sum2[696]<=1^0^Co2[695];
        Co2[696]<=(1&0|(1|0)&Co2[695]);

        Sum2[697]<=1^0^Co2[696];
        Co2[697]<=(1&0|(1|0)&Co2[696]);

        Sum2[698]<=1^0^Co2[697];
        Co2[698]<=(1&0|(1|0)&Co2[697]);

        Sum2[699]<=1^0^Co2[698];
        Co2[699]<=(1&0|(1|0)&Co2[698]);

        Sum2[700]<=1^0^Co2[699];
        Co2[700]<=(1&0|(1|0)&Co2[699]);

        Sum2[701]<=1^0^Co2[700];
        Co2[701]<=(1&0|(1|0)&Co2[700]);

        Sum2[702]<=1^0^Co2[701];
        Co2[702]<=(1&0|(1|0)&Co2[701]);

        Sum2[703]<=1^0^Co2[702];
        Co2[703]<=(1&0|(1|0)&Co2[702]);

        Sum2[704]<=1^0^Co2[703];
        Co2[704]<=(1&0|(1|0)&Co2[703]);

        Sum2[705]<=1^0^Co2[704];
        Co2[705]<=(1&0|(1|0)&Co2[704]);

        Sum2[706]<=1^0^Co2[705];
        Co2[706]<=(1&0|(1|0)&Co2[705]);

        Sum2[707]<=1^0^Co2[706];
        Co2[707]<=(1&0|(1|0)&Co2[706]);

        Sum2[708]<=1^0^Co2[707];
        Co2[708]<=(1&0|(1|0)&Co2[707]);

        Sum2[709]<=1^0^Co2[708];
        Co2[709]<=(1&0|(1|0)&Co2[708]);

        Sum2[710]<=1^0^Co2[709];
        Co2[710]<=(1&0|(1|0)&Co2[709]);

        Sum2[711]<=1^0^Co2[710];
        Co2[711]<=(1&0|(1|0)&Co2[710]);

        Sum2[712]<=1^0^Co2[711];
        Co2[712]<=(1&0|(1|0)&Co2[711]);

        Sum2[713]<=1^0^Co2[712];
        Co2[713]<=(1&0|(1|0)&Co2[712]);

        Sum2[714]<=1^0^Co2[713];
        Co2[714]<=(1&0|(1|0)&Co2[713]);

        Sum2[715]<=1^0^Co2[714];
        Co2[715]<=(1&0|(1|0)&Co2[714]);

        Sum2[716]<=1^0^Co2[715];
        Co2[716]<=(1&0|(1|0)&Co2[715]);

        Sum2[717]<=1^0^Co2[716];
        Co2[717]<=(1&0|(1|0)&Co2[716]);

        Sum2[718]<=1^0^Co2[717];
        Co2[718]<=(1&0|(1|0)&Co2[717]);

        Sum2[719]<=1^0^Co2[718];
        Co2[719]<=(1&0|(1|0)&Co2[718]);

        Sum2[720]<=1^0^Co2[719];
        Co2[720]<=(1&0|(1|0)&Co2[719]);

        Sum2[721]<=1^0^Co2[720];
        Co2[721]<=(1&0|(1|0)&Co2[720]);

        Sum2[722]<=1^0^Co2[721];
        Co2[722]<=(1&0|(1|0)&Co2[721]);

        Sum2[723]<=1^0^Co2[722];
        Co2[723]<=(1&0|(1|0)&Co2[722]);

        Sum2[724]<=1^0^Co2[723];
        Co2[724]<=(1&0|(1|0)&Co2[723]);

        Sum2[725]<=1^0^Co2[724];
        Co2[725]<=(1&0|(1|0)&Co2[724]);

        Sum2[726]<=1^0^Co2[725];
        Co2[726]<=(1&0|(1|0)&Co2[725]);

        Sum2[727]<=1^0^Co2[726];
        Co2[727]<=(1&0|(1|0)&Co2[726]);

        Sum2[728]<=1^0^Co2[727];
        Co2[728]<=(1&0|(1|0)&Co2[727]);

        Sum2[729]<=1^0^Co2[728];
        Co2[729]<=(1&0|(1|0)&Co2[728]);

        Sum2[730]<=1^0^Co2[729];
        Co2[730]<=(1&0|(1|0)&Co2[729]);

        Sum2[731]<=1^0^Co2[730];
        Co2[731]<=(1&0|(1|0)&Co2[730]);

        Sum2[732]<=1^0^Co2[731];
        Co2[732]<=(1&0|(1|0)&Co2[731]);

        Sum2[733]<=1^0^Co2[732];
        Co2[733]<=(1&0|(1|0)&Co2[732]);

        Sum2[734]<=1^0^Co2[733];
        Co2[734]<=(1&0|(1|0)&Co2[733]);

        Sum2[735]<=1^0^Co2[734];
        Co2[735]<=(1&0|(1|0)&Co2[734]);

        Sum2[736]<=1^0^Co2[735];
        Co2[736]<=(1&0|(1|0)&Co2[735]);

        Sum2[737]<=1^0^Co2[736];
        Co2[737]<=(1&0|(1|0)&Co2[736]);

        Sum2[738]<=1^0^Co2[737];
        Co2[738]<=(1&0|(1|0)&Co2[737]);

        Sum2[739]<=1^0^Co2[738];
        Co2[739]<=(1&0|(1|0)&Co2[738]);

        Sum2[740]<=1^0^Co2[739];
        Co2[740]<=(1&0|(1|0)&Co2[739]);

        Sum2[741]<=1^0^Co2[740];
        Co2[741]<=(1&0|(1|0)&Co2[740]);

        Sum2[742]<=1^0^Co2[741];
        Co2[742]<=(1&0|(1|0)&Co2[741]);

        Sum2[743]<=1^0^Co2[742];
        Co2[743]<=(1&0|(1|0)&Co2[742]);

        Sum2[744]<=1^0^Co2[743];
        Co2[744]<=(1&0|(1|0)&Co2[743]);

        Sum2[745]<=1^0^Co2[744];
        Co2[745]<=(1&0|(1|0)&Co2[744]);

        Sum2[746]<=1^0^Co2[745];
        Co2[746]<=(1&0|(1|0)&Co2[745]);

        Sum2[747]<=1^0^Co2[746];
        Co2[747]<=(1&0|(1|0)&Co2[746]);

        Sum2[748]<=1^0^Co2[747];
        Co2[748]<=(1&0|(1|0)&Co2[747]);

        Sum2[749]<=1^0^Co2[748];
        Co2[749]<=(1&0|(1|0)&Co2[748]);

        Sum2[750]<=1^0^Co2[749];
        Co2[750]<=(1&0|(1|0)&Co2[749]);

        Sum2[751]<=1^0^Co2[750];
        Co2[751]<=(1&0|(1|0)&Co2[750]);

        Sum2[752]<=1^0^Co2[751];
        Co2[752]<=(1&0|(1|0)&Co2[751]);

        Sum2[753]<=1^0^Co2[752];
        Co2[753]<=(1&0|(1|0)&Co2[752]);

        Sum2[754]<=1^0^Co2[753];
        Co2[754]<=(1&0|(1|0)&Co2[753]);

        Sum2[755]<=1^0^Co2[754];
        Co2[755]<=(1&0|(1|0)&Co2[754]);

        Sum2[756]<=1^0^Co2[755];
        Co2[756]<=(1&0|(1|0)&Co2[755]);

        Sum2[757]<=1^0^Co2[756];
        Co2[757]<=(1&0|(1|0)&Co2[756]);

        Sum2[758]<=1^0^Co2[757];
        Co2[758]<=(1&0|(1|0)&Co2[757]);

        Sum2[759]<=1^0^Co2[758];
        Co2[759]<=(1&0|(1|0)&Co2[758]);

        Sum2[760]<=1^0^Co2[759];
        Co2[760]<=(1&0|(1|0)&Co2[759]);

        Sum2[761]<=1^0^Co2[760];
        Co2[761]<=(1&0|(1|0)&Co2[760]);

        Sum2[762]<=1^0^Co2[761];
        Co2[762]<=(1&0|(1|0)&Co2[761]);

        Sum2[763]<=1^0^Co2[762];
        Co2[763]<=(1&0|(1|0)&Co2[762]);

        Sum2[764]<=1^0^Co2[763];
        Co2[764]<=(1&0|(1|0)&Co2[763]);

        Sum2[765]<=1^0^Co2[764];
        Co2[765]<=(1&0|(1|0)&Co2[764]);

        Sum2[766]<=1^0^Co2[765];
        Co2[766]<=(1&0|(1|0)&Co2[765]);

        Sum2[767]<=1^0^Co2[766];
        Co2[767]<=(1&0|(1|0)&Co2[766]);

        Sum2[768]<=1^0^Co2[767];
        Co2[768]<=(1&0|(1|0)&Co2[767]);

        Sum2[769]<=1^0^Co2[768];
        Co2[769]<=(1&0|(1|0)&Co2[768]);

        Sum2[770]<=1^0^Co2[769];
        Co2[770]<=(1&0|(1|0)&Co2[769]);

        Sum2[771]<=1^0^Co2[770];
        Co2[771]<=(1&0|(1|0)&Co2[770]);

        Sum2[772]<=1^0^Co2[771];
        Co2[772]<=(1&0|(1|0)&Co2[771]);

        Sum2[773]<=1^0^Co2[772];
        Co2[773]<=(1&0|(1|0)&Co2[772]);

        Sum2[774]<=1^0^Co2[773];
        Co2[774]<=(1&0|(1|0)&Co2[773]);

        Sum2[775]<=1^0^Co2[774];
        Co2[775]<=(1&0|(1|0)&Co2[774]);

        Sum2[776]<=1^0^Co2[775];
        Co2[776]<=(1&0|(1|0)&Co2[775]);

        Sum2[777]<=1^0^Co2[776];
        Co2[777]<=(1&0|(1|0)&Co2[776]);

        Sum2[778]<=1^0^Co2[777];
        Co2[778]<=(1&0|(1|0)&Co2[777]);

        Sum2[779]<=1^0^Co2[778];
        Co2[779]<=(1&0|(1|0)&Co2[778]);

        Sum2[780]<=1^0^Co2[779];
        Co2[780]<=(1&0|(1|0)&Co2[779]);

        Sum2[781]<=1^0^Co2[780];
        Co2[781]<=(1&0|(1|0)&Co2[780]);

        Sum2[782]<=1^0^Co2[781];
        Co2[782]<=(1&0|(1|0)&Co2[781]);

        Sum2[783]<=1^0^Co2[782];
        Co2[783]<=(1&0|(1|0)&Co2[782]);

        Sum2[784]<=1^0^Co2[783];
        Co2[784]<=(1&0|(1|0)&Co2[783]);

        Sum2[785]<=1^0^Co2[784];
        Co2[785]<=(1&0|(1|0)&Co2[784]);

        Sum2[786]<=1^0^Co2[785];
        Co2[786]<=(1&0|(1|0)&Co2[785]);

        Sum2[787]<=1^0^Co2[786];
        Co2[787]<=(1&0|(1|0)&Co2[786]);

        Sum2[788]<=1^0^Co2[787];
        Co2[788]<=(1&0|(1|0)&Co2[787]);

        Sum2[789]<=1^0^Co2[788];
        Co2[789]<=(1&0|(1|0)&Co2[788]);

        Sum2[790]<=1^0^Co2[789];
        Co2[790]<=(1&0|(1|0)&Co2[789]);

        Sum2[791]<=1^0^Co2[790];
        Co2[791]<=(1&0|(1|0)&Co2[790]);

        Sum2[792]<=1^0^Co2[791];
        Co2[792]<=(1&0|(1|0)&Co2[791]);

        Sum2[793]<=1^0^Co2[792];
        Co2[793]<=(1&0|(1|0)&Co2[792]);

        Sum2[794]<=1^0^Co2[793];
        Co2[794]<=(1&0|(1|0)&Co2[793]);

        Sum2[795]<=1^0^Co2[794];
        Co2[795]<=(1&0|(1|0)&Co2[794]);

        Sum2[796]<=1^0^Co2[795];
        Co2[796]<=(1&0|(1|0)&Co2[795]);

        Sum2[797]<=1^0^Co2[796];
        Co2[797]<=(1&0|(1|0)&Co2[796]);

        Sum2[798]<=1^0^Co2[797];
        Co2[798]<=(1&0|(1|0)&Co2[797]);

        Sum2[799]<=1^0^Co2[798];
        Co2[799]<=(1&0|(1|0)&Co2[798]);

        Sum2[800]<=1^0^Co2[799];
        Co2[800]<=(1&0|(1|0)&Co2[799]);

        Sum2[801]<=1^0^Co2[800];
        Co2[801]<=(1&0|(1|0)&Co2[800]);

        Sum2[802]<=1^0^Co2[801];
        Co2[802]<=(1&0|(1|0)&Co2[801]);

        Sum2[803]<=1^0^Co2[802];
        Co2[803]<=(1&0|(1|0)&Co2[802]);

        Sum2[804]<=1^0^Co2[803];
        Co2[804]<=(1&0|(1|0)&Co2[803]);

        Sum2[805]<=1^0^Co2[804];
        Co2[805]<=(1&0|(1|0)&Co2[804]);

        Sum2[806]<=1^0^Co2[805];
        Co2[806]<=(1&0|(1|0)&Co2[805]);

        Sum2[807]<=1^0^Co2[806];
        Co2[807]<=(1&0|(1|0)&Co2[806]);

        Sum2[808]<=1^0^Co2[807];
        Co2[808]<=(1&0|(1|0)&Co2[807]);

        Sum2[809]<=1^0^Co2[808];
        Co2[809]<=(1&0|(1|0)&Co2[808]);

        Sum2[810]<=1^0^Co2[809];
        Co2[810]<=(1&0|(1|0)&Co2[809]);

        Sum2[811]<=1^0^Co2[810];
        Co2[811]<=(1&0|(1|0)&Co2[810]);

        Sum2[812]<=1^0^Co2[811];
        Co2[812]<=(1&0|(1|0)&Co2[811]);

        Sum2[813]<=1^0^Co2[812];
        Co2[813]<=(1&0|(1|0)&Co2[812]);

        Sum2[814]<=1^0^Co2[813];
        Co2[814]<=(1&0|(1|0)&Co2[813]);

        Sum2[815]<=1^0^Co2[814];
        Co2[815]<=(1&0|(1|0)&Co2[814]);

        Sum2[816]<=1^0^Co2[815];
        Co2[816]<=(1&0|(1|0)&Co2[815]);

        Sum2[817]<=1^0^Co2[816];
        Co2[817]<=(1&0|(1|0)&Co2[816]);

        Sum2[818]<=1^0^Co2[817];
        Co2[818]<=(1&0|(1|0)&Co2[817]);

        Sum2[819]<=1^0^Co2[818];
        Co2[819]<=(1&0|(1|0)&Co2[818]);

        Sum2[820]<=1^0^Co2[819];
        Co2[820]<=(1&0|(1|0)&Co2[819]);

        Sum2[821]<=1^0^Co2[820];
        Co2[821]<=(1&0|(1|0)&Co2[820]);

        Sum2[822]<=1^0^Co2[821];
        Co2[822]<=(1&0|(1|0)&Co2[821]);

        Sum2[823]<=1^0^Co2[822];
        Co2[823]<=(1&0|(1|0)&Co2[822]);

        Sum2[824]<=1^0^Co2[823];
        Co2[824]<=(1&0|(1|0)&Co2[823]);

        Sum2[825]<=1^0^Co2[824];
        Co2[825]<=(1&0|(1|0)&Co2[824]);

        Sum2[826]<=1^0^Co2[825];
        Co2[826]<=(1&0|(1|0)&Co2[825]);

        Sum2[827]<=1^0^Co2[826];
        Co2[827]<=(1&0|(1|0)&Co2[826]);

        Sum2[828]<=1^0^Co2[827];
        Co2[828]<=(1&0|(1|0)&Co2[827]);

        Sum2[829]<=1^0^Co2[828];
        Co2[829]<=(1&0|(1|0)&Co2[828]);

        Sum2[830]<=1^0^Co2[829];
        Co2[830]<=(1&0|(1|0)&Co2[829]);

        Sum2[831]<=1^0^Co2[830];
        Co2[831]<=(1&0|(1|0)&Co2[830]);

        Sum2[832]<=1^0^Co2[831];
        Co2[832]<=(1&0|(1|0)&Co2[831]);

        Sum2[833]<=1^0^Co2[832];
        Co2[833]<=(1&0|(1|0)&Co2[832]);

        Sum2[834]<=1^0^Co2[833];
        Co2[834]<=(1&0|(1|0)&Co2[833]);

        Sum2[835]<=1^0^Co2[834];
        Co2[835]<=(1&0|(1|0)&Co2[834]);

        Sum2[836]<=1^0^Co2[835];
        Co2[836]<=(1&0|(1|0)&Co2[835]);

        Sum2[837]<=1^0^Co2[836];
        Co2[837]<=(1&0|(1|0)&Co2[836]);

        Sum2[838]<=1^0^Co2[837];
        Co2[838]<=(1&0|(1|0)&Co2[837]);

        Sum2[839]<=1^0^Co2[838];
        Co2[839]<=(1&0|(1|0)&Co2[838]);

        Sum2[840]<=1^0^Co2[839];
        Co2[840]<=(1&0|(1|0)&Co2[839]);

        Sum2[841]<=1^0^Co2[840];
        Co2[841]<=(1&0|(1|0)&Co2[840]);

        Sum2[842]<=1^0^Co2[841];
        Co2[842]<=(1&0|(1|0)&Co2[841]);

        Sum2[843]<=1^0^Co2[842];
        Co2[843]<=(1&0|(1|0)&Co2[842]);

        Sum2[844]<=1^0^Co2[843];
        Co2[844]<=(1&0|(1|0)&Co2[843]);

        Sum2[845]<=1^0^Co2[844];
        Co2[845]<=(1&0|(1|0)&Co2[844]);

        Sum2[846]<=1^0^Co2[845];
        Co2[846]<=(1&0|(1|0)&Co2[845]);

        Sum2[847]<=1^0^Co2[846];
        Co2[847]<=(1&0|(1|0)&Co2[846]);

        Sum2[848]<=1^0^Co2[847];
        Co2[848]<=(1&0|(1|0)&Co2[847]);

        Sum2[849]<=1^0^Co2[848];
        Co2[849]<=(1&0|(1|0)&Co2[848]);

        Sum2[850]<=1^0^Co2[849];
        Co2[850]<=(1&0|(1|0)&Co2[849]);

        Sum2[851]<=1^0^Co2[850];
        Co2[851]<=(1&0|(1|0)&Co2[850]);

        Sum2[852]<=1^0^Co2[851];
        Co2[852]<=(1&0|(1|0)&Co2[851]);

        Sum2[853]<=1^0^Co2[852];
        Co2[853]<=(1&0|(1|0)&Co2[852]);

        Sum2[854]<=1^0^Co2[853];
        Co2[854]<=(1&0|(1|0)&Co2[853]);

        Sum2[855]<=1^0^Co2[854];
        Co2[855]<=(1&0|(1|0)&Co2[854]);

        Sum2[856]<=1^0^Co2[855];
        Co2[856]<=(1&0|(1|0)&Co2[855]);

        Sum2[857]<=1^0^Co2[856];
        Co2[857]<=(1&0|(1|0)&Co2[856]);

        Sum2[858]<=1^0^Co2[857];
        Co2[858]<=(1&0|(1|0)&Co2[857]);

        Sum2[859]<=1^0^Co2[858];
        Co2[859]<=(1&0|(1|0)&Co2[858]);

        Sum2[860]<=1^0^Co2[859];
        Co2[860]<=(1&0|(1|0)&Co2[859]);

        Sum2[861]<=1^0^Co2[860];
        Co2[861]<=(1&0|(1|0)&Co2[860]);

        Sum2[862]<=1^0^Co2[861];
        Co2[862]<=(1&0|(1|0)&Co2[861]);

        Sum2[863]<=1^0^Co2[862];
        Co2[863]<=(1&0|(1|0)&Co2[862]);

        Sum2[864]<=1^0^Co2[863];
        Co2[864]<=(1&0|(1|0)&Co2[863]);

        Sum2[865]<=1^0^Co2[864];
        Co2[865]<=(1&0|(1|0)&Co2[864]);

        Sum2[866]<=1^0^Co2[865];
        Co2[866]<=(1&0|(1|0)&Co2[865]);

        Sum2[867]<=1^0^Co2[866];
        Co2[867]<=(1&0|(1|0)&Co2[866]);

        Sum2[868]<=1^0^Co2[867];
        Co2[868]<=(1&0|(1|0)&Co2[867]);

        Sum2[869]<=1^0^Co2[868];
        Co2[869]<=(1&0|(1|0)&Co2[868]);

        Sum2[870]<=1^0^Co2[869];
        Co2[870]<=(1&0|(1|0)&Co2[869]);

        Sum2[871]<=1^0^Co2[870];
        Co2[871]<=(1&0|(1|0)&Co2[870]);

        Sum2[872]<=1^0^Co2[871];
        Co2[872]<=(1&0|(1|0)&Co2[871]);

        Sum2[873]<=1^0^Co2[872];
        Co2[873]<=(1&0|(1|0)&Co2[872]);

        Sum2[874]<=1^0^Co2[873];
        Co2[874]<=(1&0|(1|0)&Co2[873]);

        Sum2[875]<=1^0^Co2[874];
        Co2[875]<=(1&0|(1|0)&Co2[874]);

        Sum2[876]<=1^0^Co2[875];
        Co2[876]<=(1&0|(1|0)&Co2[875]);

        Sum2[877]<=1^0^Co2[876];
        Co2[877]<=(1&0|(1|0)&Co2[876]);

        Sum2[878]<=1^0^Co2[877];
        Co2[878]<=(1&0|(1|0)&Co2[877]);

        Sum2[879]<=1^0^Co2[878];
        Co2[879]<=(1&0|(1|0)&Co2[878]);

        Sum2[880]<=1^0^Co2[879];
        Co2[880]<=(1&0|(1|0)&Co2[879]);

        Sum2[881]<=1^0^Co2[880];
        Co2[881]<=(1&0|(1|0)&Co2[880]);

        Sum2[882]<=1^0^Co2[881];
        Co2[882]<=(1&0|(1|0)&Co2[881]);

        Sum2[883]<=1^0^Co2[882];
        Co2[883]<=(1&0|(1|0)&Co2[882]);

        Sum2[884]<=1^0^Co2[883];
        Co2[884]<=(1&0|(1|0)&Co2[883]);

        Sum2[885]<=1^0^Co2[884];
        Co2[885]<=(1&0|(1|0)&Co2[884]);

        Sum2[886]<=1^0^Co2[885];
        Co2[886]<=(1&0|(1|0)&Co2[885]);

        Sum2[887]<=1^0^Co2[886];
        Co2[887]<=(1&0|(1|0)&Co2[886]);

        Sum2[888]<=1^0^Co2[887];
        Co2[888]<=(1&0|(1|0)&Co2[887]);

        Sum2[889]<=1^0^Co2[888];
        Co2[889]<=(1&0|(1|0)&Co2[888]);

        Sum2[890]<=1^0^Co2[889];
        Co2[890]<=(1&0|(1|0)&Co2[889]);

        Sum2[891]<=1^0^Co2[890];
        Co2[891]<=(1&0|(1|0)&Co2[890]);

        Sum2[892]<=1^0^Co2[891];
        Co2[892]<=(1&0|(1|0)&Co2[891]);

        Sum2[893]<=1^0^Co2[892];
        Co2[893]<=(1&0|(1|0)&Co2[892]);

        Sum2[894]<=1^0^Co2[893];
        Co2[894]<=(1&0|(1|0)&Co2[893]);

        Sum2[895]<=1^0^Co2[894];
        Co2[895]<=(1&0|(1|0)&Co2[894]);

        Sum2[896]<=1^0^Co2[895];
        Co2[896]<=(1&0|(1|0)&Co2[895]);

        Sum2[897]<=1^0^Co2[896];
        Co2[897]<=(1&0|(1|0)&Co2[896]);

        Sum2[898]<=1^0^Co2[897];
        Co2[898]<=(1&0|(1|0)&Co2[897]);

        Sum2[899]<=1^0^Co2[898];
        Co2[899]<=(1&0|(1|0)&Co2[898]);

        Sum2[900]<=1^0^Co2[899];
        Co2[900]<=(1&0|(1|0)&Co2[899]);

        Sum2[901]<=1^0^Co2[900];
        Co2[901]<=(1&0|(1|0)&Co2[900]);

        Sum2[902]<=1^0^Co2[901];
        Co2[902]<=(1&0|(1|0)&Co2[901]);

        Sum2[903]<=1^0^Co2[902];
        Co2[903]<=(1&0|(1|0)&Co2[902]);

        Sum2[904]<=1^0^Co2[903];
        Co2[904]<=(1&0|(1|0)&Co2[903]);

        Sum2[905]<=1^0^Co2[904];
        Co2[905]<=(1&0|(1|0)&Co2[904]);

        Sum2[906]<=1^0^Co2[905];
        Co2[906]<=(1&0|(1|0)&Co2[905]);

        Sum2[907]<=1^0^Co2[906];
        Co2[907]<=(1&0|(1|0)&Co2[906]);

        Sum2[908]<=1^0^Co2[907];
        Co2[908]<=(1&0|(1|0)&Co2[907]);

        Sum2[909]<=1^0^Co2[908];
        Co2[909]<=(1&0|(1|0)&Co2[908]);

        Sum2[910]<=1^0^Co2[909];
        Co2[910]<=(1&0|(1|0)&Co2[909]);

        Sum2[911]<=1^0^Co2[910];
        Co2[911]<=(1&0|(1|0)&Co2[910]);

        Sum2[912]<=1^0^Co2[911];
        Co2[912]<=(1&0|(1|0)&Co2[911]);

        Sum2[913]<=1^0^Co2[912];
        Co2[913]<=(1&0|(1|0)&Co2[912]);

        Sum2[914]<=1^0^Co2[913];
        Co2[914]<=(1&0|(1|0)&Co2[913]);

        Sum2[915]<=1^0^Co2[914];
        Co2[915]<=(1&0|(1|0)&Co2[914]);

        Sum2[916]<=1^0^Co2[915];
        Co2[916]<=(1&0|(1|0)&Co2[915]);

        Sum2[917]<=1^0^Co2[916];
        Co2[917]<=(1&0|(1|0)&Co2[916]);

        Sum2[918]<=1^0^Co2[917];
        Co2[918]<=(1&0|(1|0)&Co2[917]);

        Sum2[919]<=1^0^Co2[918];
        Co2[919]<=(1&0|(1|0)&Co2[918]);

        Sum2[920]<=1^0^Co2[919];
        Co2[920]<=(1&0|(1|0)&Co2[919]);

        Sum2[921]<=1^0^Co2[920];
        Co2[921]<=(1&0|(1|0)&Co2[920]);

        Sum2[922]<=1^0^Co2[921];
        Co2[922]<=(1&0|(1|0)&Co2[921]);

        Sum2[923]<=1^0^Co2[922];
        Co2[923]<=(1&0|(1|0)&Co2[922]);

        Sum2[924]<=1^0^Co2[923];
        Co2[924]<=(1&0|(1|0)&Co2[923]);

        Sum2[925]<=1^0^Co2[924];
        Co2[925]<=(1&0|(1|0)&Co2[924]);

        Sum2[926]<=1^0^Co2[925];
        Co2[926]<=(1&0|(1|0)&Co2[925]);

        Sum2[927]<=1^0^Co2[926];
        Co2[927]<=(1&0|(1|0)&Co2[926]);

        Sum2[928]<=1^0^Co2[927];
        Co2[928]<=(1&0|(1|0)&Co2[927]);

        Sum2[929]<=1^0^Co2[928];
        Co2[929]<=(1&0|(1|0)&Co2[928]);

        Sum2[930]<=1^0^Co2[929];
        Co2[930]<=(1&0|(1|0)&Co2[929]);

        Sum2[931]<=1^0^Co2[930];
        Co2[931]<=(1&0|(1|0)&Co2[930]);

        Sum2[932]<=1^0^Co2[931];
        Co2[932]<=(1&0|(1|0)&Co2[931]);

        Sum2[933]<=1^0^Co2[932];
        Co2[933]<=(1&0|(1|0)&Co2[932]);

        Sum2[934]<=1^0^Co2[933];
        Co2[934]<=(1&0|(1|0)&Co2[933]);

        Sum2[935]<=1^0^Co2[934];
        Co2[935]<=(1&0|(1|0)&Co2[934]);

        Sum2[936]<=1^0^Co2[935];
        Co2[936]<=(1&0|(1|0)&Co2[935]);

        Sum2[937]<=1^0^Co2[936];
        Co2[937]<=(1&0|(1|0)&Co2[936]);

        Sum2[938]<=1^0^Co2[937];
        Co2[938]<=(1&0|(1|0)&Co2[937]);

        Sum2[939]<=1^0^Co2[938];
        Co2[939]<=(1&0|(1|0)&Co2[938]);

        Sum2[940]<=1^0^Co2[939];
        Co2[940]<=(1&0|(1|0)&Co2[939]);

        Sum2[941]<=1^0^Co2[940];
        Co2[941]<=(1&0|(1|0)&Co2[940]);

        Sum2[942]<=1^0^Co2[941];
        Co2[942]<=(1&0|(1|0)&Co2[941]);

        Sum2[943]<=1^0^Co2[942];
        Co2[943]<=(1&0|(1|0)&Co2[942]);

        Sum2[944]<=1^0^Co2[943];
        Co2[944]<=(1&0|(1|0)&Co2[943]);

        Sum2[945]<=1^0^Co2[944];
        Co2[945]<=(1&0|(1|0)&Co2[944]);

        Sum2[946]<=1^0^Co2[945];
        Co2[946]<=(1&0|(1|0)&Co2[945]);

        Sum2[947]<=1^0^Co2[946];
        Co2[947]<=(1&0|(1|0)&Co2[946]);

        Sum2[948]<=1^0^Co2[947];
        Co2[948]<=(1&0|(1|0)&Co2[947]);

        Sum2[949]<=1^0^Co2[948];
        Co2[949]<=(1&0|(1|0)&Co2[948]);

        Sum2[950]<=1^0^Co2[949];
        Co2[950]<=(1&0|(1|0)&Co2[949]);

        Sum2[951]<=1^0^Co2[950];
        Co2[951]<=(1&0|(1|0)&Co2[950]);

        Sum2[952]<=1^0^Co2[951];
        Co2[952]<=(1&0|(1|0)&Co2[951]);

        Sum2[953]<=1^0^Co2[952];
        Co2[953]<=(1&0|(1|0)&Co2[952]);

        Sum2[954]<=1^0^Co2[953];
        Co2[954]<=(1&0|(1|0)&Co2[953]);

        Sum2[955]<=1^0^Co2[954];
        Co2[955]<=(1&0|(1|0)&Co2[954]);

        Sum2[956]<=1^0^Co2[955];
        Co2[956]<=(1&0|(1|0)&Co2[955]);

        Sum2[957]<=1^0^Co2[956];
        Co2[957]<=(1&0|(1|0)&Co2[956]);

        Sum2[958]<=1^0^Co2[957];
        Co2[958]<=(1&0|(1|0)&Co2[957]);

        Sum2[959]<=1^0^Co2[958];
        Co2[959]<=(1&0|(1|0)&Co2[958]);

        Sum2[960]<=1^0^Co2[959];
        Co2[960]<=(1&0|(1|0)&Co2[959]);

        Sum2[961]<=1^0^Co2[960];
        Co2[961]<=(1&0|(1|0)&Co2[960]);

        Sum2[962]<=1^0^Co2[961];
        Co2[962]<=(1&0|(1|0)&Co2[961]);

        Sum2[963]<=1^0^Co2[962];
        Co2[963]<=(1&0|(1|0)&Co2[962]);

        Sum2[964]<=1^0^Co2[963];
        Co2[964]<=(1&0|(1|0)&Co2[963]);

        Sum2[965]<=1^0^Co2[964];
        Co2[965]<=(1&0|(1|0)&Co2[964]);

        Sum2[966]<=1^0^Co2[965];
        Co2[966]<=(1&0|(1|0)&Co2[965]);

        Sum2[967]<=1^0^Co2[966];
        Co2[967]<=(1&0|(1|0)&Co2[966]);

        Sum2[968]<=1^0^Co2[967];
        Co2[968]<=(1&0|(1|0)&Co2[967]);

        Sum2[969]<=1^0^Co2[968];
        Co2[969]<=(1&0|(1|0)&Co2[968]);

        Sum2[970]<=1^0^Co2[969];
        Co2[970]<=(1&0|(1|0)&Co2[969]);

        Sum2[971]<=1^0^Co2[970];
        Co2[971]<=(1&0|(1|0)&Co2[970]);

        Sum2[972]<=1^0^Co2[971];
        Co2[972]<=(1&0|(1|0)&Co2[971]);

        Sum2[973]<=1^0^Co2[972];
        Co2[973]<=(1&0|(1|0)&Co2[972]);

        Sum2[974]<=1^0^Co2[973];
        Co2[974]<=(1&0|(1|0)&Co2[973]);

        Sum2[975]<=1^0^Co2[974];
        Co2[975]<=(1&0|(1|0)&Co2[974]);

        Sum2[976]<=1^0^Co2[975];
        Co2[976]<=(1&0|(1|0)&Co2[975]);

        Sum2[977]<=1^0^Co2[976];
        Co2[977]<=(1&0|(1|0)&Co2[976]);

        Sum2[978]<=1^0^Co2[977];
        Co2[978]<=(1&0|(1|0)&Co2[977]);

        Sum2[979]<=1^0^Co2[978];
        Co2[979]<=(1&0|(1|0)&Co2[978]);

        Sum2[980]<=1^0^Co2[979];
        Co2[980]<=(1&0|(1|0)&Co2[979]);

        Sum2[981]<=1^0^Co2[980];
        Co2[981]<=(1&0|(1|0)&Co2[980]);

        Sum2[982]<=1^0^Co2[981];
        Co2[982]<=(1&0|(1|0)&Co2[981]);

        Sum2[983]<=1^0^Co2[982];
        Co2[983]<=(1&0|(1|0)&Co2[982]);

        Sum2[984]<=1^0^Co2[983];
        Co2[984]<=(1&0|(1|0)&Co2[983]);

        Sum2[985]<=1^0^Co2[984];
        Co2[985]<=(1&0|(1|0)&Co2[984]);

        Sum2[986]<=1^0^Co2[985];
        Co2[986]<=(1&0|(1|0)&Co2[985]);

        Sum2[987]<=1^0^Co2[986];
        Co2[987]<=(1&0|(1|0)&Co2[986]);

        Sum2[988]<=1^0^Co2[987];
        Co2[988]<=(1&0|(1|0)&Co2[987]);

        Sum2[989]<=1^0^Co2[988];
        Co2[989]<=(1&0|(1|0)&Co2[988]);

        Sum2[990]<=1^0^Co2[989];
        Co2[990]<=(1&0|(1|0)&Co2[989]);

        Sum2[991]<=1^0^Co2[990];
        Co2[991]<=(1&0|(1|0)&Co2[990]);

        Sum2[992]<=1^0^Co2[991];
        Co2[992]<=(1&0|(1|0)&Co2[991]);

        Sum2[993]<=1^0^Co2[992];
        Co2[993]<=(1&0|(1|0)&Co2[992]);

        Sum2[994]<=1^0^Co2[993];
        Co2[994]<=(1&0|(1|0)&Co2[993]);

        Sum2[995]<=1^0^Co2[994];
        Co2[995]<=(1&0|(1|0)&Co2[994]);

        Sum2[996]<=1^0^Co2[995];
        Co2[996]<=(1&0|(1|0)&Co2[995]);

        Sum2[997]<=1^0^Co2[996];
        Co2[997]<=(1&0|(1|0)&Co2[996]);

        Sum2[998]<=1^0^Co2[997];
        Co2[998]<=(1&0|(1|0)&Co2[997]);

        Sum2[999]<=1^0^Co2[998];
        Co2[999]<=(1&0|(1|0)&Co2[998]);

        Sum2[1000]<=1^0^Co2[999];
        Co2[1000]<=(1&0|(1|0)&Co2[999]);

        Sum2[1001]<=1^0^Co2[1000];
        Co2[1001]<=(1&0|(1|0)&Co2[1000]);

        Sum2[1002]<=1^0^Co2[1001];
        Co2[1002]<=(1&0|(1|0)&Co2[1001]);

        Sum2[1003]<=1^0^Co2[1002];
        Co2[1003]<=(1&0|(1|0)&Co2[1002]);

        Sum2[1004]<=1^0^Co2[1003];
        Co2[1004]<=(1&0|(1|0)&Co2[1003]);

        Sum2[1005]<=1^0^Co2[1004];
        Co2[1005]<=(1&0|(1|0)&Co2[1004]);

        Sum2[1006]<=1^0^Co2[1005];
        Co2[1006]<=(1&0|(1|0)&Co2[1005]);

        Sum2[1007]<=1^0^Co2[1006];
        Co2[1007]<=(1&0|(1|0)&Co2[1006]);

        Sum2[1008]<=1^0^Co2[1007];
        Co2[1008]<=(1&0|(1|0)&Co2[1007]);

        Sum2[1009]<=1^0^Co2[1008];
        Co2[1009]<=(1&0|(1|0)&Co2[1008]);

        Sum2[1010]<=1^0^Co2[1009];
        Co2[1010]<=(1&0|(1|0)&Co2[1009]);

        Sum2[1011]<=1^0^Co2[1010];
        Co2[1011]<=(1&0|(1|0)&Co2[1010]);

        Sum2[1012]<=1^0^Co2[1011];
        Co2[1012]<=(1&0|(1|0)&Co2[1011]);

        Sum2[1013]<=1^0^Co2[1012];
        Co2[1013]<=(1&0|(1|0)&Co2[1012]);

        Sum2[1014]<=1^0^Co2[1013];
        Co2[1014]<=(1&0|(1|0)&Co2[1013]);

        Sum2[1015]<=1^0^Co2[1014];
        Co2[1015]<=(1&0|(1|0)&Co2[1014]);

        Sum2[1016]<=1^0^Co2[1015];
        Co2[1016]<=(1&0|(1|0)&Co2[1015]);

        Sum2[1017]<=1^0^Co2[1016];
        Co2[1017]<=(1&0|(1|0)&Co2[1016]);

        Sum2[1018]<=1^0^Co2[1017];
        Co2[1018]<=(1&0|(1|0)&Co2[1017]);

        Sum2[1019]<=1^0^Co2[1018];
        Co2[1019]<=(1&0|(1|0)&Co2[1018]);

        Sum2[1020]<=1^0^Co2[1019];
        Co2[1020]<=(1&0|(1|0)&Co2[1019]);

        Sum2[1021]<=1^0^Co2[1020];
        Co2[1021]<=(1&0|(1|0)&Co2[1020]);

        Sum2[1022]<=1^0^Co2[1021];
        Co2[1022]<=(1&0|(1|0)&Co2[1021]);

        Sum2[1023]<=1^0^Co2[1022];
        Co2[1023]<=(1&0|(1|0)&Co2[1022]);

        // part 2
        /*
        LED1 <= 1;
        Sum2[1023:0] <= 4096'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
        Co2[1023:0] <= 4096'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
                Sum2[0]<=1^Hit^Ci;
        Co2[0]<=(1&Hit|(1|Hit)&Ci);

        Sum2[1]<=1^0^Co2[0];
        Co2[1]<=(1&0|(1|0)&Co2[0]);

        Sum2[2]<=1^0^Co2[1];
        Co2[2]<=(1&0|(1|0)&Co2[1]);

        Sum2[3]<=1^0^Co2[2];
        Co2[3]<=(1&0|(1|0)&Co2[2]);

        Sum2[4]<=1^0^Co2[3];
        Co2[4]<=(1&0|(1|0)&Co2[3]);

        Sum2[5]<=1^0^Co2[4];
        Co2[5]<=(1&0|(1|0)&Co2[4]);

        Sum2[6]<=1^0^Co2[5];
        Co2[6]<=(1&0|(1|0)&Co2[5]);

        Sum2[7]<=1^0^Co2[6];
        Co2[7]<=(1&0|(1|0)&Co2[6]);

        Sum2[8]<=1^0^Co2[7];
        Co2[8]<=(1&0|(1|0)&Co2[7]);

        Sum2[9]<=1^0^Co2[8];
        Co2[9]<=(1&0|(1|0)&Co2[8]);

        Sum2[10]<=1^0^Co2[9];
        Co2[10]<=(1&0|(1|0)&Co2[9]);

        Sum2[11]<=1^0^Co2[10];
        Co2[11]<=(1&0|(1|0)&Co2[10]);

        Sum2[12]<=1^0^Co2[11];
        Co2[12]<=(1&0|(1|0)&Co2[11]);

        Sum2[13]<=1^0^Co2[12];
        Co2[13]<=(1&0|(1|0)&Co2[12]);

        Sum2[14]<=1^0^Co2[13];
        Co2[14]<=(1&0|(1|0)&Co2[13]);

        Sum2[15]<=1^0^Co2[14];
        Co2[15]<=(1&0|(1|0)&Co2[14]);

        Sum2[16]<=1^0^Co2[15];
        Co2[16]<=(1&0|(1|0)&Co2[15]);

        Sum2[17]<=1^0^Co2[16];
        Co2[17]<=(1&0|(1|0)&Co2[16]);

        Sum2[18]<=1^0^Co2[17];
        Co2[18]<=(1&0|(1|0)&Co2[17]);

        Sum2[19]<=1^0^Co2[18];
        Co2[19]<=(1&0|(1|0)&Co2[18]);

        Sum2[20]<=1^0^Co2[19];
        Co2[20]<=(1&0|(1|0)&Co2[19]);

        Sum2[21]<=1^0^Co2[20];
        Co2[21]<=(1&0|(1|0)&Co2[20]);

        Sum2[22]<=1^0^Co2[21];
        Co2[22]<=(1&0|(1|0)&Co2[21]);

        Sum2[23]<=1^0^Co2[22];
        Co2[23]<=(1&0|(1|0)&Co2[22]);

        Sum2[24]<=1^0^Co2[23];
        Co2[24]<=(1&0|(1|0)&Co2[23]);

        Sum2[25]<=1^0^Co2[24];
        Co2[25]<=(1&0|(1|0)&Co2[24]);

        Sum2[26]<=1^0^Co2[25];
        Co2[26]<=(1&0|(1|0)&Co2[25]);

        Sum2[27]<=1^0^Co2[26];
        Co2[27]<=(1&0|(1|0)&Co2[26]);

        Sum2[28]<=1^0^Co2[27];
        Co2[28]<=(1&0|(1|0)&Co2[27]);

        Sum2[29]<=1^0^Co2[28];
        Co2[29]<=(1&0|(1|0)&Co2[28]);

        Sum2[30]<=1^0^Co2[29];
        Co2[30]<=(1&0|(1|0)&Co2[29]);

        Sum2[31]<=1^0^Co2[30];
        Co2[31]<=(1&0|(1|0)&Co2[30]);

        Sum2[32]<=1^0^Co2[31];
        Co2[32]<=(1&0|(1|0)&Co2[31]);

        Sum2[33]<=1^0^Co2[32];
        Co2[33]<=(1&0|(1|0)&Co2[32]);

        Sum2[34]<=1^0^Co2[33];
        Co2[34]<=(1&0|(1|0)&Co2[33]);

        Sum2[35]<=1^0^Co2[34];
        Co2[35]<=(1&0|(1|0)&Co2[34]);

        Sum2[36]<=1^0^Co2[35];
        Co2[36]<=(1&0|(1|0)&Co2[35]);

        Sum2[37]<=1^0^Co2[36];
        Co2[37]<=(1&0|(1|0)&Co2[36]);

        Sum2[38]<=1^0^Co2[37];
        Co2[38]<=(1&0|(1|0)&Co2[37]);

        Sum2[39]<=1^0^Co2[38];
        Co2[39]<=(1&0|(1|0)&Co2[38]);

        Sum2[40]<=1^0^Co2[39];
        Co2[40]<=(1&0|(1|0)&Co2[39]);

        Sum2[41]<=1^0^Co2[40];
        Co2[41]<=(1&0|(1|0)&Co2[40]);

        Sum2[42]<=1^0^Co2[41];
        Co2[42]<=(1&0|(1|0)&Co2[41]);

        Sum2[43]<=1^0^Co2[42];
        Co2[43]<=(1&0|(1|0)&Co2[42]);

        Sum2[44]<=1^0^Co2[43];
        Co2[44]<=(1&0|(1|0)&Co2[43]);

        Sum2[45]<=1^0^Co2[44];
        Co2[45]<=(1&0|(1|0)&Co2[44]);

        Sum2[46]<=1^0^Co2[45];
        Co2[46]<=(1&0|(1|0)&Co2[45]);

        Sum2[47]<=1^0^Co2[46];
        Co2[47]<=(1&0|(1|0)&Co2[46]);

        Sum2[48]<=1^0^Co2[47];
        Co2[48]<=(1&0|(1|0)&Co2[47]);

        Sum2[49]<=1^0^Co2[48];
        Co2[49]<=(1&0|(1|0)&Co2[48]);

        Sum2[50]<=1^0^Co2[49];
        Co2[50]<=(1&0|(1|0)&Co2[49]);

        Sum2[51]<=1^0^Co2[50];
        Co2[51]<=(1&0|(1|0)&Co2[50]);

        Sum2[52]<=1^0^Co2[51];
        Co2[52]<=(1&0|(1|0)&Co2[51]);

        Sum2[53]<=1^0^Co2[52];
        Co2[53]<=(1&0|(1|0)&Co2[52]);

        Sum2[54]<=1^0^Co2[53];
        Co2[54]<=(1&0|(1|0)&Co2[53]);

        Sum2[55]<=1^0^Co2[54];
        Co2[55]<=(1&0|(1|0)&Co2[54]);

        Sum2[56]<=1^0^Co2[55];
        Co2[56]<=(1&0|(1|0)&Co2[55]);

        Sum2[57]<=1^0^Co2[56];
        Co2[57]<=(1&0|(1|0)&Co2[56]);

        Sum2[58]<=1^0^Co2[57];
        Co2[58]<=(1&0|(1|0)&Co2[57]);

        Sum2[59]<=1^0^Co2[58];
        Co2[59]<=(1&0|(1|0)&Co2[58]);

        Sum2[60]<=1^0^Co2[59];
        Co2[60]<=(1&0|(1|0)&Co2[59]);

        Sum2[61]<=1^0^Co2[60];
        Co2[61]<=(1&0|(1|0)&Co2[60]);

        Sum2[62]<=1^0^Co2[61];
        Co2[62]<=(1&0|(1|0)&Co2[61]);

        Sum2[63]<=1^0^Co2[62];
        Co2[63]<=(1&0|(1|0)&Co2[62]);

        Sum2[64]<=1^0^Co2[63];
        Co2[64]<=(1&0|(1|0)&Co2[63]);

        Sum2[65]<=1^0^Co2[64];
        Co2[65]<=(1&0|(1|0)&Co2[64]);

        Sum2[66]<=1^0^Co2[65];
        Co2[66]<=(1&0|(1|0)&Co2[65]);

        Sum2[67]<=1^0^Co2[66];
        Co2[67]<=(1&0|(1|0)&Co2[66]);

        Sum2[68]<=1^0^Co2[67];
        Co2[68]<=(1&0|(1|0)&Co2[67]);

        Sum2[69]<=1^0^Co2[68];
        Co2[69]<=(1&0|(1|0)&Co2[68]);

        Sum2[70]<=1^0^Co2[69];
        Co2[70]<=(1&0|(1|0)&Co2[69]);

        Sum2[71]<=1^0^Co2[70];
        Co2[71]<=(1&0|(1|0)&Co2[70]);

        Sum2[72]<=1^0^Co2[71];
        Co2[72]<=(1&0|(1|0)&Co2[71]);

        Sum2[73]<=1^0^Co2[72];
        Co2[73]<=(1&0|(1|0)&Co2[72]);

        Sum2[74]<=1^0^Co2[73];
        Co2[74]<=(1&0|(1|0)&Co2[73]);

        Sum2[75]<=1^0^Co2[74];
        Co2[75]<=(1&0|(1|0)&Co2[74]);

        Sum2[76]<=1^0^Co2[75];
        Co2[76]<=(1&0|(1|0)&Co2[75]);

        Sum2[77]<=1^0^Co2[76];
        Co2[77]<=(1&0|(1|0)&Co2[76]);

        Sum2[78]<=1^0^Co2[77];
        Co2[78]<=(1&0|(1|0)&Co2[77]);

        Sum2[79]<=1^0^Co2[78];
        Co2[79]<=(1&0|(1|0)&Co2[78]);

        Sum2[80]<=1^0^Co2[79];
        Co2[80]<=(1&0|(1|0)&Co2[79]);

        Sum2[81]<=1^0^Co2[80];
        Co2[81]<=(1&0|(1|0)&Co2[80]);

        Sum2[82]<=1^0^Co2[81];
        Co2[82]<=(1&0|(1|0)&Co2[81]);

        Sum2[83]<=1^0^Co2[82];
        Co2[83]<=(1&0|(1|0)&Co2[82]);

        Sum2[84]<=1^0^Co2[83];
        Co2[84]<=(1&0|(1|0)&Co2[83]);

        Sum2[85]<=1^0^Co2[84];
        Co2[85]<=(1&0|(1|0)&Co2[84]);

        Sum2[86]<=1^0^Co2[85];
        Co2[86]<=(1&0|(1|0)&Co2[85]);

        Sum2[87]<=1^0^Co2[86];
        Co2[87]<=(1&0|(1|0)&Co2[86]);

        Sum2[88]<=1^0^Co2[87];
        Co2[88]<=(1&0|(1|0)&Co2[87]);

        Sum2[89]<=1^0^Co2[88];
        Co2[89]<=(1&0|(1|0)&Co2[88]);

        Sum2[90]<=1^0^Co2[89];
        Co2[90]<=(1&0|(1|0)&Co2[89]);

        Sum2[91]<=1^0^Co2[90];
        Co2[91]<=(1&0|(1|0)&Co2[90]);

        Sum2[92]<=1^0^Co2[91];
        Co2[92]<=(1&0|(1|0)&Co2[91]);

        Sum2[93]<=1^0^Co2[92];
        Co2[93]<=(1&0|(1|0)&Co2[92]);

        Sum2[94]<=1^0^Co2[93];
        Co2[94]<=(1&0|(1|0)&Co2[93]);

        Sum2[95]<=1^0^Co2[94];
        Co2[95]<=(1&0|(1|0)&Co2[94]);

        Sum2[96]<=1^0^Co2[95];
        Co2[96]<=(1&0|(1|0)&Co2[95]);

        Sum2[97]<=1^0^Co2[96];
        Co2[97]<=(1&0|(1|0)&Co2[96]);

        Sum2[98]<=1^0^Co2[97];
        Co2[98]<=(1&0|(1|0)&Co2[97]);

        Sum2[99]<=1^0^Co2[98];
        Co2[99]<=(1&0|(1|0)&Co2[98]);

        Sum2[100]<=1^0^Co2[99];
        Co2[100]<=(1&0|(1|0)&Co2[99]);

        Sum2[101]<=1^0^Co2[100];
        Co2[101]<=(1&0|(1|0)&Co2[100]);

        Sum2[102]<=1^0^Co2[101];
        Co2[102]<=(1&0|(1|0)&Co2[101]);

        Sum2[103]<=1^0^Co2[102];
        Co2[103]<=(1&0|(1|0)&Co2[102]);

        Sum2[104]<=1^0^Co2[103];
        Co2[104]<=(1&0|(1|0)&Co2[103]);

        Sum2[105]<=1^0^Co2[104];
        Co2[105]<=(1&0|(1|0)&Co2[104]);

        Sum2[106]<=1^0^Co2[105];
        Co2[106]<=(1&0|(1|0)&Co2[105]);

        Sum2[107]<=1^0^Co2[106];
        Co2[107]<=(1&0|(1|0)&Co2[106]);

        Sum2[108]<=1^0^Co2[107];
        Co2[108]<=(1&0|(1|0)&Co2[107]);

        Sum2[109]<=1^0^Co2[108];
        Co2[109]<=(1&0|(1|0)&Co2[108]);

        Sum2[110]<=1^0^Co2[109];
        Co2[110]<=(1&0|(1|0)&Co2[109]);

        Sum2[111]<=1^0^Co2[110];
        Co2[111]<=(1&0|(1|0)&Co2[110]);

        Sum2[112]<=1^0^Co2[111];
        Co2[112]<=(1&0|(1|0)&Co2[111]);

        Sum2[113]<=1^0^Co2[112];
        Co2[113]<=(1&0|(1|0)&Co2[112]);

        Sum2[114]<=1^0^Co2[113];
        Co2[114]<=(1&0|(1|0)&Co2[113]);

        Sum2[115]<=1^0^Co2[114];
        Co2[115]<=(1&0|(1|0)&Co2[114]);

        Sum2[116]<=1^0^Co2[115];
        Co2[116]<=(1&0|(1|0)&Co2[115]);

        Sum2[117]<=1^0^Co2[116];
        Co2[117]<=(1&0|(1|0)&Co2[116]);

        Sum2[118]<=1^0^Co2[117];
        Co2[118]<=(1&0|(1|0)&Co2[117]);

        Sum2[119]<=1^0^Co2[118];
        Co2[119]<=(1&0|(1|0)&Co2[118]);

        Sum2[120]<=1^0^Co2[119];
        Co2[120]<=(1&0|(1|0)&Co2[119]);

        Sum2[121]<=1^0^Co2[120];
        Co2[121]<=(1&0|(1|0)&Co2[120]);

        Sum2[122]<=1^0^Co2[121];
        Co2[122]<=(1&0|(1|0)&Co2[121]);

        Sum2[123]<=1^0^Co2[122];
        Co2[123]<=(1&0|(1|0)&Co2[122]);

        Sum2[124]<=1^0^Co2[123];
        Co2[124]<=(1&0|(1|0)&Co2[123]);

        Sum2[125]<=1^0^Co2[124];
        Co2[125]<=(1&0|(1|0)&Co2[124]);

        Sum2[126]<=1^0^Co2[125];
        Co2[126]<=(1&0|(1|0)&Co2[125]);

        Sum2[127]<=1^0^Co2[126];
        Co2[127]<=(1&0|(1|0)&Co2[126]);

        Sum2[128]<=1^0^Co2[127];
        Co2[128]<=(1&0|(1|0)&Co2[127]);

        Sum2[129]<=1^0^Co2[128];
        Co2[129]<=(1&0|(1|0)&Co2[128]);

        Sum2[130]<=1^0^Co2[129];
        Co2[130]<=(1&0|(1|0)&Co2[129]);

        Sum2[131]<=1^0^Co2[130];
        Co2[131]<=(1&0|(1|0)&Co2[130]);

        Sum2[132]<=1^0^Co2[131];
        Co2[132]<=(1&0|(1|0)&Co2[131]);

        Sum2[133]<=1^0^Co2[132];
        Co2[133]<=(1&0|(1|0)&Co2[132]);

        Sum2[134]<=1^0^Co2[133];
        Co2[134]<=(1&0|(1|0)&Co2[133]);

        Sum2[135]<=1^0^Co2[134];
        Co2[135]<=(1&0|(1|0)&Co2[134]);

        Sum2[136]<=1^0^Co2[135];
        Co2[136]<=(1&0|(1|0)&Co2[135]);

        Sum2[137]<=1^0^Co2[136];
        Co2[137]<=(1&0|(1|0)&Co2[136]);

        Sum2[138]<=1^0^Co2[137];
        Co2[138]<=(1&0|(1|0)&Co2[137]);

        Sum2[139]<=1^0^Co2[138];
        Co2[139]<=(1&0|(1|0)&Co2[138]);

        Sum2[140]<=1^0^Co2[139];
        Co2[140]<=(1&0|(1|0)&Co2[139]);

        Sum2[141]<=1^0^Co2[140];
        Co2[141]<=(1&0|(1|0)&Co2[140]);

        Sum2[142]<=1^0^Co2[141];
        Co2[142]<=(1&0|(1|0)&Co2[141]);

        Sum2[143]<=1^0^Co2[142];
        Co2[143]<=(1&0|(1|0)&Co2[142]);

        Sum2[144]<=1^0^Co2[143];
        Co2[144]<=(1&0|(1|0)&Co2[143]);

        Sum2[145]<=1^0^Co2[144];
        Co2[145]<=(1&0|(1|0)&Co2[144]);

        Sum2[146]<=1^0^Co2[145];
        Co2[146]<=(1&0|(1|0)&Co2[145]);

        Sum2[147]<=1^0^Co2[146];
        Co2[147]<=(1&0|(1|0)&Co2[146]);

        Sum2[148]<=1^0^Co2[147];
        Co2[148]<=(1&0|(1|0)&Co2[147]);

        Sum2[149]<=1^0^Co2[148];
        Co2[149]<=(1&0|(1|0)&Co2[148]);

        Sum2[150]<=1^0^Co2[149];
        Co2[150]<=(1&0|(1|0)&Co2[149]);

        Sum2[151]<=1^0^Co2[150];
        Co2[151]<=(1&0|(1|0)&Co2[150]);

        Sum2[152]<=1^0^Co2[151];
        Co2[152]<=(1&0|(1|0)&Co2[151]);

        Sum2[153]<=1^0^Co2[152];
        Co2[153]<=(1&0|(1|0)&Co2[152]);

        Sum2[154]<=1^0^Co2[153];
        Co2[154]<=(1&0|(1|0)&Co2[153]);

        Sum2[155]<=1^0^Co2[154];
        Co2[155]<=(1&0|(1|0)&Co2[154]);

        Sum2[156]<=1^0^Co2[155];
        Co2[156]<=(1&0|(1|0)&Co2[155]);

        Sum2[157]<=1^0^Co2[156];
        Co2[157]<=(1&0|(1|0)&Co2[156]);

        Sum2[158]<=1^0^Co2[157];
        Co2[158]<=(1&0|(1|0)&Co2[157]);

        Sum2[159]<=1^0^Co2[158];
        Co2[159]<=(1&0|(1|0)&Co2[158]);

        Sum2[160]<=1^0^Co2[159];
        Co2[160]<=(1&0|(1|0)&Co2[159]);

        Sum2[161]<=1^0^Co2[160];
        Co2[161]<=(1&0|(1|0)&Co2[160]);

        Sum2[162]<=1^0^Co2[161];
        Co2[162]<=(1&0|(1|0)&Co2[161]);

        Sum2[163]<=1^0^Co2[162];
        Co2[163]<=(1&0|(1|0)&Co2[162]);

        Sum2[164]<=1^0^Co2[163];
        Co2[164]<=(1&0|(1|0)&Co2[163]);

        Sum2[165]<=1^0^Co2[164];
        Co2[165]<=(1&0|(1|0)&Co2[164]);

        Sum2[166]<=1^0^Co2[165];
        Co2[166]<=(1&0|(1|0)&Co2[165]);

        Sum2[167]<=1^0^Co2[166];
        Co2[167]<=(1&0|(1|0)&Co2[166]);

        Sum2[168]<=1^0^Co2[167];
        Co2[168]<=(1&0|(1|0)&Co2[167]);

        Sum2[169]<=1^0^Co2[168];
        Co2[169]<=(1&0|(1|0)&Co2[168]);

        Sum2[170]<=1^0^Co2[169];
        Co2[170]<=(1&0|(1|0)&Co2[169]);

        Sum2[171]<=1^0^Co2[170];
        Co2[171]<=(1&0|(1|0)&Co2[170]);

        Sum2[172]<=1^0^Co2[171];
        Co2[172]<=(1&0|(1|0)&Co2[171]);

        Sum2[173]<=1^0^Co2[172];
        Co2[173]<=(1&0|(1|0)&Co2[172]);

        Sum2[174]<=1^0^Co2[173];
        Co2[174]<=(1&0|(1|0)&Co2[173]);

        Sum2[175]<=1^0^Co2[174];
        Co2[175]<=(1&0|(1|0)&Co2[174]);

        Sum2[176]<=1^0^Co2[175];
        Co2[176]<=(1&0|(1|0)&Co2[175]);

        Sum2[177]<=1^0^Co2[176];
        Co2[177]<=(1&0|(1|0)&Co2[176]);

        Sum2[178]<=1^0^Co2[177];
        Co2[178]<=(1&0|(1|0)&Co2[177]);

        Sum2[179]<=1^0^Co2[178];
        Co2[179]<=(1&0|(1|0)&Co2[178]);

        Sum2[180]<=1^0^Co2[179];
        Co2[180]<=(1&0|(1|0)&Co2[179]);

        Sum2[181]<=1^0^Co2[180];
        Co2[181]<=(1&0|(1|0)&Co2[180]);

        Sum2[182]<=1^0^Co2[181];
        Co2[182]<=(1&0|(1|0)&Co2[181]);

        Sum2[183]<=1^0^Co2[182];
        Co2[183]<=(1&0|(1|0)&Co2[182]);

        Sum2[184]<=1^0^Co2[183];
        Co2[184]<=(1&0|(1|0)&Co2[183]);

        Sum2[185]<=1^0^Co2[184];
        Co2[185]<=(1&0|(1|0)&Co2[184]);

        Sum2[186]<=1^0^Co2[185];
        Co2[186]<=(1&0|(1|0)&Co2[185]);

        Sum2[187]<=1^0^Co2[186];
        Co2[187]<=(1&0|(1|0)&Co2[186]);

        Sum2[188]<=1^0^Co2[187];
        Co2[188]<=(1&0|(1|0)&Co2[187]);

        Sum2[189]<=1^0^Co2[188];
        Co2[189]<=(1&0|(1|0)&Co2[188]);

        Sum2[190]<=1^0^Co2[189];
        Co2[190]<=(1&0|(1|0)&Co2[189]);

        Sum2[191]<=1^0^Co2[190];
        Co2[191]<=(1&0|(1|0)&Co2[190]);

        Sum2[192]<=1^0^Co2[191];
        Co2[192]<=(1&0|(1|0)&Co2[191]);

        Sum2[193]<=1^0^Co2[192];
        Co2[193]<=(1&0|(1|0)&Co2[192]);

        Sum2[194]<=1^0^Co2[193];
        Co2[194]<=(1&0|(1|0)&Co2[193]);

        Sum2[195]<=1^0^Co2[194];
        Co2[195]<=(1&0|(1|0)&Co2[194]);

        Sum2[196]<=1^0^Co2[195];
        Co2[196]<=(1&0|(1|0)&Co2[195]);

        Sum2[197]<=1^0^Co2[196];
        Co2[197]<=(1&0|(1|0)&Co2[196]);

        Sum2[198]<=1^0^Co2[197];
        Co2[198]<=(1&0|(1|0)&Co2[197]);

        Sum2[199]<=1^0^Co2[198];
        Co2[199]<=(1&0|(1|0)&Co2[198]);

        Sum2[200]<=1^0^Co2[199];
        Co2[200]<=(1&0|(1|0)&Co2[199]);

        Sum2[201]<=1^0^Co2[200];
        Co2[201]<=(1&0|(1|0)&Co2[200]);

        Sum2[202]<=1^0^Co2[201];
        Co2[202]<=(1&0|(1|0)&Co2[201]);

        Sum2[203]<=1^0^Co2[202];
        Co2[203]<=(1&0|(1|0)&Co2[202]);

        Sum2[204]<=1^0^Co2[203];
        Co2[204]<=(1&0|(1|0)&Co2[203]);

        Sum2[205]<=1^0^Co2[204];
        Co2[205]<=(1&0|(1|0)&Co2[204]);

        Sum2[206]<=1^0^Co2[205];
        Co2[206]<=(1&0|(1|0)&Co2[205]);

        Sum2[207]<=1^0^Co2[206];
        Co2[207]<=(1&0|(1|0)&Co2[206]);

        Sum2[208]<=1^0^Co2[207];
        Co2[208]<=(1&0|(1|0)&Co2[207]);

        Sum2[209]<=1^0^Co2[208];
        Co2[209]<=(1&0|(1|0)&Co2[208]);

        Sum2[210]<=1^0^Co2[209];
        Co2[210]<=(1&0|(1|0)&Co2[209]);

        Sum2[211]<=1^0^Co2[210];
        Co2[211]<=(1&0|(1|0)&Co2[210]);

        Sum2[212]<=1^0^Co2[211];
        Co2[212]<=(1&0|(1|0)&Co2[211]);

        Sum2[213]<=1^0^Co2[212];
        Co2[213]<=(1&0|(1|0)&Co2[212]);

        Sum2[214]<=1^0^Co2[213];
        Co2[214]<=(1&0|(1|0)&Co2[213]);

        Sum2[215]<=1^0^Co2[214];
        Co2[215]<=(1&0|(1|0)&Co2[214]);

        Sum2[216]<=1^0^Co2[215];
        Co2[216]<=(1&0|(1|0)&Co2[215]);

        Sum2[217]<=1^0^Co2[216];
        Co2[217]<=(1&0|(1|0)&Co2[216]);

        Sum2[218]<=1^0^Co2[217];
        Co2[218]<=(1&0|(1|0)&Co2[217]);

        Sum2[219]<=1^0^Co2[218];
        Co2[219]<=(1&0|(1|0)&Co2[218]);

        Sum2[220]<=1^0^Co2[219];
        Co2[220]<=(1&0|(1|0)&Co2[219]);

        Sum2[221]<=1^0^Co2[220];
        Co2[221]<=(1&0|(1|0)&Co2[220]);

        Sum2[222]<=1^0^Co2[221];
        Co2[222]<=(1&0|(1|0)&Co2[221]);

        Sum2[223]<=1^0^Co2[222];
        Co2[223]<=(1&0|(1|0)&Co2[222]);

        Sum2[224]<=1^0^Co2[223];
        Co2[224]<=(1&0|(1|0)&Co2[223]);

        Sum2[225]<=1^0^Co2[224];
        Co2[225]<=(1&0|(1|0)&Co2[224]);

        Sum2[226]<=1^0^Co2[225];
        Co2[226]<=(1&0|(1|0)&Co2[225]);

        Sum2[227]<=1^0^Co2[226];
        Co2[227]<=(1&0|(1|0)&Co2[226]);

        Sum2[228]<=1^0^Co2[227];
        Co2[228]<=(1&0|(1|0)&Co2[227]);

        Sum2[229]<=1^0^Co2[228];
        Co2[229]<=(1&0|(1|0)&Co2[228]);

        Sum2[230]<=1^0^Co2[229];
        Co2[230]<=(1&0|(1|0)&Co2[229]);

        Sum2[231]<=1^0^Co2[230];
        Co2[231]<=(1&0|(1|0)&Co2[230]);

        Sum2[232]<=1^0^Co2[231];
        Co2[232]<=(1&0|(1|0)&Co2[231]);

        Sum2[233]<=1^0^Co2[232];
        Co2[233]<=(1&0|(1|0)&Co2[232]);

        Sum2[234]<=1^0^Co2[233];
        Co2[234]<=(1&0|(1|0)&Co2[233]);

        Sum2[235]<=1^0^Co2[234];
        Co2[235]<=(1&0|(1|0)&Co2[234]);

        Sum2[236]<=1^0^Co2[235];
        Co2[236]<=(1&0|(1|0)&Co2[235]);

        Sum2[237]<=1^0^Co2[236];
        Co2[237]<=(1&0|(1|0)&Co2[236]);

        Sum2[238]<=1^0^Co2[237];
        Co2[238]<=(1&0|(1|0)&Co2[237]);

        Sum2[239]<=1^0^Co2[238];
        Co2[239]<=(1&0|(1|0)&Co2[238]);

        Sum2[240]<=1^0^Co2[239];
        Co2[240]<=(1&0|(1|0)&Co2[239]);

        Sum2[241]<=1^0^Co2[240];
        Co2[241]<=(1&0|(1|0)&Co2[240]);

        Sum2[242]<=1^0^Co2[241];
        Co2[242]<=(1&0|(1|0)&Co2[241]);

        Sum2[243]<=1^0^Co2[242];
        Co2[243]<=(1&0|(1|0)&Co2[242]);

        Sum2[244]<=1^0^Co2[243];
        Co2[244]<=(1&0|(1|0)&Co2[243]);

        Sum2[245]<=1^0^Co2[244];
        Co2[245]<=(1&0|(1|0)&Co2[244]);

        Sum2[246]<=1^0^Co2[245];
        Co2[246]<=(1&0|(1|0)&Co2[245]);

        Sum2[247]<=1^0^Co2[246];
        Co2[247]<=(1&0|(1|0)&Co2[246]);

        Sum2[248]<=1^0^Co2[247];
        Co2[248]<=(1&0|(1|0)&Co2[247]);

        Sum2[249]<=1^0^Co2[248];
        Co2[249]<=(1&0|(1|0)&Co2[248]);

        Sum2[250]<=1^0^Co2[249];
        Co2[250]<=(1&0|(1|0)&Co2[249]);

        Sum2[251]<=1^0^Co2[250];
        Co2[251]<=(1&0|(1|0)&Co2[250]);

        Sum2[252]<=1^0^Co2[251];
        Co2[252]<=(1&0|(1|0)&Co2[251]);

        Sum2[253]<=1^0^Co2[252];
        Co2[253]<=(1&0|(1|0)&Co2[252]);

        Sum2[254]<=1^0^Co2[253];
        Co2[254]<=(1&0|(1|0)&Co2[253]);

        Sum2[255]<=1^0^Co2[254];
        Co2[255]<=(1&0|(1|0)&Co2[254]);

        Sum2[256]<=1^0^Co2[255];
        Co2[256]<=(1&0|(1|0)&Co2[255]);

        Sum2[257]<=1^0^Co2[256];
        Co2[257]<=(1&0|(1|0)&Co2[256]);

        Sum2[258]<=1^0^Co2[257];
        Co2[258]<=(1&0|(1|0)&Co2[257]);

        Sum2[259]<=1^0^Co2[258];
        Co2[259]<=(1&0|(1|0)&Co2[258]);

        Sum2[260]<=1^0^Co2[259];
        Co2[260]<=(1&0|(1|0)&Co2[259]);

        Sum2[261]<=1^0^Co2[260];
        Co2[261]<=(1&0|(1|0)&Co2[260]);

        Sum2[262]<=1^0^Co2[261];
        Co2[262]<=(1&0|(1|0)&Co2[261]);

        Sum2[263]<=1^0^Co2[262];
        Co2[263]<=(1&0|(1|0)&Co2[262]);

        Sum2[264]<=1^0^Co2[263];
        Co2[264]<=(1&0|(1|0)&Co2[263]);

        Sum2[265]<=1^0^Co2[264];
        Co2[265]<=(1&0|(1|0)&Co2[264]);

        Sum2[266]<=1^0^Co2[265];
        Co2[266]<=(1&0|(1|0)&Co2[265]);

        Sum2[267]<=1^0^Co2[266];
        Co2[267]<=(1&0|(1|0)&Co2[266]);

        Sum2[268]<=1^0^Co2[267];
        Co2[268]<=(1&0|(1|0)&Co2[267]);

        Sum2[269]<=1^0^Co2[268];
        Co2[269]<=(1&0|(1|0)&Co2[268]);

        Sum2[270]<=1^0^Co2[269];
        Co2[270]<=(1&0|(1|0)&Co2[269]);

        Sum2[271]<=1^0^Co2[270];
        Co2[271]<=(1&0|(1|0)&Co2[270]);

        Sum2[272]<=1^0^Co2[271];
        Co2[272]<=(1&0|(1|0)&Co2[271]);

        Sum2[273]<=1^0^Co2[272];
        Co2[273]<=(1&0|(1|0)&Co2[272]);

        Sum2[274]<=1^0^Co2[273];
        Co2[274]<=(1&0|(1|0)&Co2[273]);

        Sum2[275]<=1^0^Co2[274];
        Co2[275]<=(1&0|(1|0)&Co2[274]);

        Sum2[276]<=1^0^Co2[275];
        Co2[276]<=(1&0|(1|0)&Co2[275]);

        Sum2[277]<=1^0^Co2[276];
        Co2[277]<=(1&0|(1|0)&Co2[276]);

        Sum2[278]<=1^0^Co2[277];
        Co2[278]<=(1&0|(1|0)&Co2[277]);

        Sum2[279]<=1^0^Co2[278];
        Co2[279]<=(1&0|(1|0)&Co2[278]);

        Sum2[280]<=1^0^Co2[279];
        Co2[280]<=(1&0|(1|0)&Co2[279]);

        Sum2[281]<=1^0^Co2[280];
        Co2[281]<=(1&0|(1|0)&Co2[280]);

        Sum2[282]<=1^0^Co2[281];
        Co2[282]<=(1&0|(1|0)&Co2[281]);

        Sum2[283]<=1^0^Co2[282];
        Co2[283]<=(1&0|(1|0)&Co2[282]);

        Sum2[284]<=1^0^Co2[283];
        Co2[284]<=(1&0|(1|0)&Co2[283]);

        Sum2[285]<=1^0^Co2[284];
        Co2[285]<=(1&0|(1|0)&Co2[284]);

        Sum2[286]<=1^0^Co2[285];
        Co2[286]<=(1&0|(1|0)&Co2[285]);

        Sum2[287]<=1^0^Co2[286];
        Co2[287]<=(1&0|(1|0)&Co2[286]);

        Sum2[288]<=1^0^Co2[287];
        Co2[288]<=(1&0|(1|0)&Co2[287]);

        Sum2[289]<=1^0^Co2[288];
        Co2[289]<=(1&0|(1|0)&Co2[288]);

        Sum2[290]<=1^0^Co2[289];
        Co2[290]<=(1&0|(1|0)&Co2[289]);

        Sum2[291]<=1^0^Co2[290];
        Co2[291]<=(1&0|(1|0)&Co2[290]);

        Sum2[292]<=1^0^Co2[291];
        Co2[292]<=(1&0|(1|0)&Co2[291]);

        Sum2[293]<=1^0^Co2[292];
        Co2[293]<=(1&0|(1|0)&Co2[292]);

        Sum2[294]<=1^0^Co2[293];
        Co2[294]<=(1&0|(1|0)&Co2[293]);

        Sum2[295]<=1^0^Co2[294];
        Co2[295]<=(1&0|(1|0)&Co2[294]);

        Sum2[296]<=1^0^Co2[295];
        Co2[296]<=(1&0|(1|0)&Co2[295]);

        Sum2[297]<=1^0^Co2[296];
        Co2[297]<=(1&0|(1|0)&Co2[296]);

        Sum2[298]<=1^0^Co2[297];
        Co2[298]<=(1&0|(1|0)&Co2[297]);

        Sum2[299]<=1^0^Co2[298];
        Co2[299]<=(1&0|(1|0)&Co2[298]);

        Sum2[300]<=1^0^Co2[299];
        Co2[300]<=(1&0|(1|0)&Co2[299]);

        Sum2[301]<=1^0^Co2[300];
        Co2[301]<=(1&0|(1|0)&Co2[300]);

        Sum2[302]<=1^0^Co2[301];
        Co2[302]<=(1&0|(1|0)&Co2[301]);

        Sum2[303]<=1^0^Co2[302];
        Co2[303]<=(1&0|(1|0)&Co2[302]);

        Sum2[304]<=1^0^Co2[303];
        Co2[304]<=(1&0|(1|0)&Co2[303]);

        Sum2[305]<=1^0^Co2[304];
        Co2[305]<=(1&0|(1|0)&Co2[304]);

        Sum2[306]<=1^0^Co2[305];
        Co2[306]<=(1&0|(1|0)&Co2[305]);

        Sum2[307]<=1^0^Co2[306];
        Co2[307]<=(1&0|(1|0)&Co2[306]);

        Sum2[308]<=1^0^Co2[307];
        Co2[308]<=(1&0|(1|0)&Co2[307]);

        Sum2[309]<=1^0^Co2[308];
        Co2[309]<=(1&0|(1|0)&Co2[308]);

        Sum2[310]<=1^0^Co2[309];
        Co2[310]<=(1&0|(1|0)&Co2[309]);

        Sum2[311]<=1^0^Co2[310];
        Co2[311]<=(1&0|(1|0)&Co2[310]);

        Sum2[312]<=1^0^Co2[311];
        Co2[312]<=(1&0|(1|0)&Co2[311]);

        Sum2[313]<=1^0^Co2[312];
        Co2[313]<=(1&0|(1|0)&Co2[312]);

        Sum2[314]<=1^0^Co2[313];
        Co2[314]<=(1&0|(1|0)&Co2[313]);

        Sum2[315]<=1^0^Co2[314];
        Co2[315]<=(1&0|(1|0)&Co2[314]);

        Sum2[316]<=1^0^Co2[315];
        Co2[316]<=(1&0|(1|0)&Co2[315]);

        Sum2[317]<=1^0^Co2[316];
        Co2[317]<=(1&0|(1|0)&Co2[316]);

        Sum2[318]<=1^0^Co2[317];
        Co2[318]<=(1&0|(1|0)&Co2[317]);

        Sum2[319]<=1^0^Co2[318];
        Co2[319]<=(1&0|(1|0)&Co2[318]);

        Sum2[320]<=1^0^Co2[319];
        Co2[320]<=(1&0|(1|0)&Co2[319]);

        Sum2[321]<=1^0^Co2[320];
        Co2[321]<=(1&0|(1|0)&Co2[320]);

        Sum2[322]<=1^0^Co2[321];
        Co2[322]<=(1&0|(1|0)&Co2[321]);

        Sum2[323]<=1^0^Co2[322];
        Co2[323]<=(1&0|(1|0)&Co2[322]);

        Sum2[324]<=1^0^Co2[323];
        Co2[324]<=(1&0|(1|0)&Co2[323]);

        Sum2[325]<=1^0^Co2[324];
        Co2[325]<=(1&0|(1|0)&Co2[324]);

        Sum2[326]<=1^0^Co2[325];
        Co2[326]<=(1&0|(1|0)&Co2[325]);

        Sum2[327]<=1^0^Co2[326];
        Co2[327]<=(1&0|(1|0)&Co2[326]);

        Sum2[328]<=1^0^Co2[327];
        Co2[328]<=(1&0|(1|0)&Co2[327]);

        Sum2[329]<=1^0^Co2[328];
        Co2[329]<=(1&0|(1|0)&Co2[328]);

        Sum2[330]<=1^0^Co2[329];
        Co2[330]<=(1&0|(1|0)&Co2[329]);

        Sum2[331]<=1^0^Co2[330];
        Co2[331]<=(1&0|(1|0)&Co2[330]);

        Sum2[332]<=1^0^Co2[331];
        Co2[332]<=(1&0|(1|0)&Co2[331]);

        Sum2[333]<=1^0^Co2[332];
        Co2[333]<=(1&0|(1|0)&Co2[332]);

        Sum2[334]<=1^0^Co2[333];
        Co2[334]<=(1&0|(1|0)&Co2[333]);

        Sum2[335]<=1^0^Co2[334];
        Co2[335]<=(1&0|(1|0)&Co2[334]);

        Sum2[336]<=1^0^Co2[335];
        Co2[336]<=(1&0|(1|0)&Co2[335]);

        Sum2[337]<=1^0^Co2[336];
        Co2[337]<=(1&0|(1|0)&Co2[336]);

        Sum2[338]<=1^0^Co2[337];
        Co2[338]<=(1&0|(1|0)&Co2[337]);

        Sum2[339]<=1^0^Co2[338];
        Co2[339]<=(1&0|(1|0)&Co2[338]);

        Sum2[340]<=1^0^Co2[339];
        Co2[340]<=(1&0|(1|0)&Co2[339]);

        Sum2[341]<=1^0^Co2[340];
        Co2[341]<=(1&0|(1|0)&Co2[340]);

        Sum2[342]<=1^0^Co2[341];
        Co2[342]<=(1&0|(1|0)&Co2[341]);

        Sum2[343]<=1^0^Co2[342];
        Co2[343]<=(1&0|(1|0)&Co2[342]);

        Sum2[344]<=1^0^Co2[343];
        Co2[344]<=(1&0|(1|0)&Co2[343]);

        Sum2[345]<=1^0^Co2[344];
        Co2[345]<=(1&0|(1|0)&Co2[344]);

        Sum2[346]<=1^0^Co2[345];
        Co2[346]<=(1&0|(1|0)&Co2[345]);

        Sum2[347]<=1^0^Co2[346];
        Co2[347]<=(1&0|(1|0)&Co2[346]);

        Sum2[348]<=1^0^Co2[347];
        Co2[348]<=(1&0|(1|0)&Co2[347]);

        Sum2[349]<=1^0^Co2[348];
        Co2[349]<=(1&0|(1|0)&Co2[348]);

        Sum2[350]<=1^0^Co2[349];
        Co2[350]<=(1&0|(1|0)&Co2[349]);

        Sum2[351]<=1^0^Co2[350];
        Co2[351]<=(1&0|(1|0)&Co2[350]);

        Sum2[352]<=1^0^Co2[351];
        Co2[352]<=(1&0|(1|0)&Co2[351]);

        Sum2[353]<=1^0^Co2[352];
        Co2[353]<=(1&0|(1|0)&Co2[352]);

        Sum2[354]<=1^0^Co2[353];
        Co2[354]<=(1&0|(1|0)&Co2[353]);

        Sum2[355]<=1^0^Co2[354];
        Co2[355]<=(1&0|(1|0)&Co2[354]);

        Sum2[356]<=1^0^Co2[355];
        Co2[356]<=(1&0|(1|0)&Co2[355]);

        Sum2[357]<=1^0^Co2[356];
        Co2[357]<=(1&0|(1|0)&Co2[356]);

        Sum2[358]<=1^0^Co2[357];
        Co2[358]<=(1&0|(1|0)&Co2[357]);

        Sum2[359]<=1^0^Co2[358];
        Co2[359]<=(1&0|(1|0)&Co2[358]);

        Sum2[360]<=1^0^Co2[359];
        Co2[360]<=(1&0|(1|0)&Co2[359]);

        Sum2[361]<=1^0^Co2[360];
        Co2[361]<=(1&0|(1|0)&Co2[360]);

        Sum2[362]<=1^0^Co2[361];
        Co2[362]<=(1&0|(1|0)&Co2[361]);

        Sum2[363]<=1^0^Co2[362];
        Co2[363]<=(1&0|(1|0)&Co2[362]);

        Sum2[364]<=1^0^Co2[363];
        Co2[364]<=(1&0|(1|0)&Co2[363]);

        Sum2[365]<=1^0^Co2[364];
        Co2[365]<=(1&0|(1|0)&Co2[364]);

        Sum2[366]<=1^0^Co2[365];
        Co2[366]<=(1&0|(1|0)&Co2[365]);

        Sum2[367]<=1^0^Co2[366];
        Co2[367]<=(1&0|(1|0)&Co2[366]);

        Sum2[368]<=1^0^Co2[367];
        Co2[368]<=(1&0|(1|0)&Co2[367]);

        Sum2[369]<=1^0^Co2[368];
        Co2[369]<=(1&0|(1|0)&Co2[368]);

        Sum2[370]<=1^0^Co2[369];
        Co2[370]<=(1&0|(1|0)&Co2[369]);

        Sum2[371]<=1^0^Co2[370];
        Co2[371]<=(1&0|(1|0)&Co2[370]);

        Sum2[372]<=1^0^Co2[371];
        Co2[372]<=(1&0|(1|0)&Co2[371]);

        Sum2[373]<=1^0^Co2[372];
        Co2[373]<=(1&0|(1|0)&Co2[372]);

        Sum2[374]<=1^0^Co2[373];
        Co2[374]<=(1&0|(1|0)&Co2[373]);

        Sum2[375]<=1^0^Co2[374];
        Co2[375]<=(1&0|(1|0)&Co2[374]);

        Sum2[376]<=1^0^Co2[375];
        Co2[376]<=(1&0|(1|0)&Co2[375]);

        Sum2[377]<=1^0^Co2[376];
        Co2[377]<=(1&0|(1|0)&Co2[376]);

        Sum2[378]<=1^0^Co2[377];
        Co2[378]<=(1&0|(1|0)&Co2[377]);

        Sum2[379]<=1^0^Co2[378];
        Co2[379]<=(1&0|(1|0)&Co2[378]);

        Sum2[380]<=1^0^Co2[379];
        Co2[380]<=(1&0|(1|0)&Co2[379]);

        Sum2[381]<=1^0^Co2[380];
        Co2[381]<=(1&0|(1|0)&Co2[380]);

        Sum2[382]<=1^0^Co2[381];
        Co2[382]<=(1&0|(1|0)&Co2[381]);

        Sum2[383]<=1^0^Co2[382];
        Co2[383]<=(1&0|(1|0)&Co2[382]);

        Sum2[384]<=1^0^Co2[383];
        Co2[384]<=(1&0|(1|0)&Co2[383]);

        Sum2[385]<=1^0^Co2[384];
        Co2[385]<=(1&0|(1|0)&Co2[384]);

        Sum2[386]<=1^0^Co2[385];
        Co2[386]<=(1&0|(1|0)&Co2[385]);

        Sum2[387]<=1^0^Co2[386];
        Co2[387]<=(1&0|(1|0)&Co2[386]);

        Sum2[388]<=1^0^Co2[387];
        Co2[388]<=(1&0|(1|0)&Co2[387]);

        Sum2[389]<=1^0^Co2[388];
        Co2[389]<=(1&0|(1|0)&Co2[388]);

        Sum2[390]<=1^0^Co2[389];
        Co2[390]<=(1&0|(1|0)&Co2[389]);

        Sum2[391]<=1^0^Co2[390];
        Co2[391]<=(1&0|(1|0)&Co2[390]);

        Sum2[392]<=1^0^Co2[391];
        Co2[392]<=(1&0|(1|0)&Co2[391]);

        Sum2[393]<=1^0^Co2[392];
        Co2[393]<=(1&0|(1|0)&Co2[392]);

        Sum2[394]<=1^0^Co2[393];
        Co2[394]<=(1&0|(1|0)&Co2[393]);

        Sum2[395]<=1^0^Co2[394];
        Co2[395]<=(1&0|(1|0)&Co2[394]);

        Sum2[396]<=1^0^Co2[395];
        Co2[396]<=(1&0|(1|0)&Co2[395]);

        Sum2[397]<=1^0^Co2[396];
        Co2[397]<=(1&0|(1|0)&Co2[396]);

        Sum2[398]<=1^0^Co2[397];
        Co2[398]<=(1&0|(1|0)&Co2[397]);

        Sum2[399]<=1^0^Co2[398];
        Co2[399]<=(1&0|(1|0)&Co2[398]);

        Sum2[400]<=1^0^Co2[399];
        Co2[400]<=(1&0|(1|0)&Co2[399]);

        Sum2[401]<=1^0^Co2[400];
        Co2[401]<=(1&0|(1|0)&Co2[400]);

        Sum2[402]<=1^0^Co2[401];
        Co2[402]<=(1&0|(1|0)&Co2[401]);

        Sum2[403]<=1^0^Co2[402];
        Co2[403]<=(1&0|(1|0)&Co2[402]);

        Sum2[404]<=1^0^Co2[403];
        Co2[404]<=(1&0|(1|0)&Co2[403]);

        Sum2[405]<=1^0^Co2[404];
        Co2[405]<=(1&0|(1|0)&Co2[404]);

        Sum2[406]<=1^0^Co2[405];
        Co2[406]<=(1&0|(1|0)&Co2[405]);

        Sum2[407]<=1^0^Co2[406];
        Co2[407]<=(1&0|(1|0)&Co2[406]);

        Sum2[408]<=1^0^Co2[407];
        Co2[408]<=(1&0|(1|0)&Co2[407]);

        Sum2[409]<=1^0^Co2[408];
        Co2[409]<=(1&0|(1|0)&Co2[408]);

        Sum2[410]<=1^0^Co2[409];
        Co2[410]<=(1&0|(1|0)&Co2[409]);

        Sum2[411]<=1^0^Co2[410];
        Co2[411]<=(1&0|(1|0)&Co2[410]);

        Sum2[412]<=1^0^Co2[411];
        Co2[412]<=(1&0|(1|0)&Co2[411]);

        Sum2[413]<=1^0^Co2[412];
        Co2[413]<=(1&0|(1|0)&Co2[412]);

        Sum2[414]<=1^0^Co2[413];
        Co2[414]<=(1&0|(1|0)&Co2[413]);

        Sum2[415]<=1^0^Co2[414];
        Co2[415]<=(1&0|(1|0)&Co2[414]);

        Sum2[416]<=1^0^Co2[415];
        Co2[416]<=(1&0|(1|0)&Co2[415]);

        Sum2[417]<=1^0^Co2[416];
        Co2[417]<=(1&0|(1|0)&Co2[416]);

        Sum2[418]<=1^0^Co2[417];
        Co2[418]<=(1&0|(1|0)&Co2[417]);

        Sum2[419]<=1^0^Co2[418];
        Co2[419]<=(1&0|(1|0)&Co2[418]);

        Sum2[420]<=1^0^Co2[419];
        Co2[420]<=(1&0|(1|0)&Co2[419]);

        Sum2[421]<=1^0^Co2[420];
        Co2[421]<=(1&0|(1|0)&Co2[420]);

        Sum2[422]<=1^0^Co2[421];
        Co2[422]<=(1&0|(1|0)&Co2[421]);

        Sum2[423]<=1^0^Co2[422];
        Co2[423]<=(1&0|(1|0)&Co2[422]);

        Sum2[424]<=1^0^Co2[423];
        Co2[424]<=(1&0|(1|0)&Co2[423]);

        Sum2[425]<=1^0^Co2[424];
        Co2[425]<=(1&0|(1|0)&Co2[424]);

        Sum2[426]<=1^0^Co2[425];
        Co2[426]<=(1&0|(1|0)&Co2[425]);

        Sum2[427]<=1^0^Co2[426];
        Co2[427]<=(1&0|(1|0)&Co2[426]);

        Sum2[428]<=1^0^Co2[427];
        Co2[428]<=(1&0|(1|0)&Co2[427]);

        Sum2[429]<=1^0^Co2[428];
        Co2[429]<=(1&0|(1|0)&Co2[428]);

        Sum2[430]<=1^0^Co2[429];
        Co2[430]<=(1&0|(1|0)&Co2[429]);

        Sum2[431]<=1^0^Co2[430];
        Co2[431]<=(1&0|(1|0)&Co2[430]);

        Sum2[432]<=1^0^Co2[431];
        Co2[432]<=(1&0|(1|0)&Co2[431]);

        Sum2[433]<=1^0^Co2[432];
        Co2[433]<=(1&0|(1|0)&Co2[432]);

        Sum2[434]<=1^0^Co2[433];
        Co2[434]<=(1&0|(1|0)&Co2[433]);

        Sum2[435]<=1^0^Co2[434];
        Co2[435]<=(1&0|(1|0)&Co2[434]);

        Sum2[436]<=1^0^Co2[435];
        Co2[436]<=(1&0|(1|0)&Co2[435]);

        Sum2[437]<=1^0^Co2[436];
        Co2[437]<=(1&0|(1|0)&Co2[436]);

        Sum2[438]<=1^0^Co2[437];
        Co2[438]<=(1&0|(1|0)&Co2[437]);

        Sum2[439]<=1^0^Co2[438];
        Co2[439]<=(1&0|(1|0)&Co2[438]);

        Sum2[440]<=1^0^Co2[439];
        Co2[440]<=(1&0|(1|0)&Co2[439]);

        Sum2[441]<=1^0^Co2[440];
        Co2[441]<=(1&0|(1|0)&Co2[440]);

        Sum2[442]<=1^0^Co2[441];
        Co2[442]<=(1&0|(1|0)&Co2[441]);

        Sum2[443]<=1^0^Co2[442];
        Co2[443]<=(1&0|(1|0)&Co2[442]);

        Sum2[444]<=1^0^Co2[443];
        Co2[444]<=(1&0|(1|0)&Co2[443]);

        Sum2[445]<=1^0^Co2[444];
        Co2[445]<=(1&0|(1|0)&Co2[444]);

        Sum2[446]<=1^0^Co2[445];
        Co2[446]<=(1&0|(1|0)&Co2[445]);

        Sum2[447]<=1^0^Co2[446];
        Co2[447]<=(1&0|(1|0)&Co2[446]);

        Sum2[448]<=1^0^Co2[447];
        Co2[448]<=(1&0|(1|0)&Co2[447]);

        Sum2[449]<=1^0^Co2[448];
        Co2[449]<=(1&0|(1|0)&Co2[448]);

        Sum2[450]<=1^0^Co2[449];
        Co2[450]<=(1&0|(1|0)&Co2[449]);

        Sum2[451]<=1^0^Co2[450];
        Co2[451]<=(1&0|(1|0)&Co2[450]);

        Sum2[452]<=1^0^Co2[451];
        Co2[452]<=(1&0|(1|0)&Co2[451]);

        Sum2[453]<=1^0^Co2[452];
        Co2[453]<=(1&0|(1|0)&Co2[452]);

        Sum2[454]<=1^0^Co2[453];
        Co2[454]<=(1&0|(1|0)&Co2[453]);

        Sum2[455]<=1^0^Co2[454];
        Co2[455]<=(1&0|(1|0)&Co2[454]);

        Sum2[456]<=1^0^Co2[455];
        Co2[456]<=(1&0|(1|0)&Co2[455]);

        Sum2[457]<=1^0^Co2[456];
        Co2[457]<=(1&0|(1|0)&Co2[456]);

        Sum2[458]<=1^0^Co2[457];
        Co2[458]<=(1&0|(1|0)&Co2[457]);

        Sum2[459]<=1^0^Co2[458];
        Co2[459]<=(1&0|(1|0)&Co2[458]);

        Sum2[460]<=1^0^Co2[459];
        Co2[460]<=(1&0|(1|0)&Co2[459]);

        Sum2[461]<=1^0^Co2[460];
        Co2[461]<=(1&0|(1|0)&Co2[460]);

        Sum2[462]<=1^0^Co2[461];
        Co2[462]<=(1&0|(1|0)&Co2[461]);

        Sum2[463]<=1^0^Co2[462];
        Co2[463]<=(1&0|(1|0)&Co2[462]);

        Sum2[464]<=1^0^Co2[463];
        Co2[464]<=(1&0|(1|0)&Co2[463]);

        Sum2[465]<=1^0^Co2[464];
        Co2[465]<=(1&0|(1|0)&Co2[464]);

        Sum2[466]<=1^0^Co2[465];
        Co2[466]<=(1&0|(1|0)&Co2[465]);

        Sum2[467]<=1^0^Co2[466];
        Co2[467]<=(1&0|(1|0)&Co2[466]);

        Sum2[468]<=1^0^Co2[467];
        Co2[468]<=(1&0|(1|0)&Co2[467]);

        Sum2[469]<=1^0^Co2[468];
        Co2[469]<=(1&0|(1|0)&Co2[468]);

        Sum2[470]<=1^0^Co2[469];
        Co2[470]<=(1&0|(1|0)&Co2[469]);

        Sum2[471]<=1^0^Co2[470];
        Co2[471]<=(1&0|(1|0)&Co2[470]);

        Sum2[472]<=1^0^Co2[471];
        Co2[472]<=(1&0|(1|0)&Co2[471]);

        Sum2[473]<=1^0^Co2[472];
        Co2[473]<=(1&0|(1|0)&Co2[472]);

        Sum2[474]<=1^0^Co2[473];
        Co2[474]<=(1&0|(1|0)&Co2[473]);

        Sum2[475]<=1^0^Co2[474];
        Co2[475]<=(1&0|(1|0)&Co2[474]);

        Sum2[476]<=1^0^Co2[475];
        Co2[476]<=(1&0|(1|0)&Co2[475]);

        Sum2[477]<=1^0^Co2[476];
        Co2[477]<=(1&0|(1|0)&Co2[476]);

        Sum2[478]<=1^0^Co2[477];
        Co2[478]<=(1&0|(1|0)&Co2[477]);

        Sum2[479]<=1^0^Co2[478];
        Co2[479]<=(1&0|(1|0)&Co2[478]);

        Sum2[480]<=1^0^Co2[479];
        Co2[480]<=(1&0|(1|0)&Co2[479]);

        Sum2[481]<=1^0^Co2[480];
        Co2[481]<=(1&0|(1|0)&Co2[480]);

        Sum2[482]<=1^0^Co2[481];
        Co2[482]<=(1&0|(1|0)&Co2[481]);

        Sum2[483]<=1^0^Co2[482];
        Co2[483]<=(1&0|(1|0)&Co2[482]);

        Sum2[484]<=1^0^Co2[483];
        Co2[484]<=(1&0|(1|0)&Co2[483]);

        Sum2[485]<=1^0^Co2[484];
        Co2[485]<=(1&0|(1|0)&Co2[484]);

        Sum2[486]<=1^0^Co2[485];
        Co2[486]<=(1&0|(1|0)&Co2[485]);

        Sum2[487]<=1^0^Co2[486];
        Co2[487]<=(1&0|(1|0)&Co2[486]);

        Sum2[488]<=1^0^Co2[487];
        Co2[488]<=(1&0|(1|0)&Co2[487]);

        Sum2[489]<=1^0^Co2[488];
        Co2[489]<=(1&0|(1|0)&Co2[488]);

        Sum2[490]<=1^0^Co2[489];
        Co2[490]<=(1&0|(1|0)&Co2[489]);

        Sum2[491]<=1^0^Co2[490];
        Co2[491]<=(1&0|(1|0)&Co2[490]);

        Sum2[492]<=1^0^Co2[491];
        Co2[492]<=(1&0|(1|0)&Co2[491]);

        Sum2[493]<=1^0^Co2[492];
        Co2[493]<=(1&0|(1|0)&Co2[492]);

        Sum2[494]<=1^0^Co2[493];
        Co2[494]<=(1&0|(1|0)&Co2[493]);

        Sum2[495]<=1^0^Co2[494];
        Co2[495]<=(1&0|(1|0)&Co2[494]);

        Sum2[496]<=1^0^Co2[495];
        Co2[496]<=(1&0|(1|0)&Co2[495]);

        Sum2[497]<=1^0^Co2[496];
        Co2[497]<=(1&0|(1|0)&Co2[496]);

        Sum2[498]<=1^0^Co2[497];
        Co2[498]<=(1&0|(1|0)&Co2[497]);

        Sum2[499]<=1^0^Co2[498];
        Co2[499]<=(1&0|(1|0)&Co2[498]);

        Sum2[500]<=1^0^Co2[499];
        Co2[500]<=(1&0|(1|0)&Co2[499]);

        Sum2[501]<=1^0^Co2[500];
        Co2[501]<=(1&0|(1|0)&Co2[500]);

        Sum2[502]<=1^0^Co2[501];
        Co2[502]<=(1&0|(1|0)&Co2[501]);

        Sum2[503]<=1^0^Co2[502];
        Co2[503]<=(1&0|(1|0)&Co2[502]);

        Sum2[504]<=1^0^Co2[503];
        Co2[504]<=(1&0|(1|0)&Co2[503]);

        Sum2[505]<=1^0^Co2[504];
        Co2[505]<=(1&0|(1|0)&Co2[504]);

        Sum2[506]<=1^0^Co2[505];
        Co2[506]<=(1&0|(1|0)&Co2[505]);

        Sum2[507]<=1^0^Co2[506];
        Co2[507]<=(1&0|(1|0)&Co2[506]);

        Sum2[508]<=1^0^Co2[507];
        Co2[508]<=(1&0|(1|0)&Co2[507]);

        Sum2[509]<=1^0^Co2[508];
        Co2[509]<=(1&0|(1|0)&Co2[508]);

        Sum2[510]<=1^0^Co2[509];
        Co2[510]<=(1&0|(1|0)&Co2[509]);

        Sum2[511]<=1^0^Co2[510];
        Co2[511]<=(1&0|(1|0)&Co2[510]);

        Sum2[512]<=1^0^Co2[511];
        Co2[512]<=(1&0|(1|0)&Co2[511]);

        Sum2[513]<=1^0^Co2[512];
        Co2[513]<=(1&0|(1|0)&Co2[512]);

        Sum2[514]<=1^0^Co2[513];
        Co2[514]<=(1&0|(1|0)&Co2[513]);

        Sum2[515]<=1^0^Co2[514];
        Co2[515]<=(1&0|(1|0)&Co2[514]);

        Sum2[516]<=1^0^Co2[515];
        Co2[516]<=(1&0|(1|0)&Co2[515]);

        Sum2[517]<=1^0^Co2[516];
        Co2[517]<=(1&0|(1|0)&Co2[516]);

        Sum2[518]<=1^0^Co2[517];
        Co2[518]<=(1&0|(1|0)&Co2[517]);

        Sum2[519]<=1^0^Co2[518];
        Co2[519]<=(1&0|(1|0)&Co2[518]);

        Sum2[520]<=1^0^Co2[519];
        Co2[520]<=(1&0|(1|0)&Co2[519]);

        Sum2[521]<=1^0^Co2[520];
        Co2[521]<=(1&0|(1|0)&Co2[520]);

        Sum2[522]<=1^0^Co2[521];
        Co2[522]<=(1&0|(1|0)&Co2[521]);

        Sum2[523]<=1^0^Co2[522];
        Co2[523]<=(1&0|(1|0)&Co2[522]);

        Sum2[524]<=1^0^Co2[523];
        Co2[524]<=(1&0|(1|0)&Co2[523]);

        Sum2[525]<=1^0^Co2[524];
        Co2[525]<=(1&0|(1|0)&Co2[524]);

        Sum2[526]<=1^0^Co2[525];
        Co2[526]<=(1&0|(1|0)&Co2[525]);

        Sum2[527]<=1^0^Co2[526];
        Co2[527]<=(1&0|(1|0)&Co2[526]);

        Sum2[528]<=1^0^Co2[527];
        Co2[528]<=(1&0|(1|0)&Co2[527]);

        Sum2[529]<=1^0^Co2[528];
        Co2[529]<=(1&0|(1|0)&Co2[528]);

        Sum2[530]<=1^0^Co2[529];
        Co2[530]<=(1&0|(1|0)&Co2[529]);

        Sum2[531]<=1^0^Co2[530];
        Co2[531]<=(1&0|(1|0)&Co2[530]);

        Sum2[532]<=1^0^Co2[531];
        Co2[532]<=(1&0|(1|0)&Co2[531]);

        Sum2[533]<=1^0^Co2[532];
        Co2[533]<=(1&0|(1|0)&Co2[532]);

        Sum2[534]<=1^0^Co2[533];
        Co2[534]<=(1&0|(1|0)&Co2[533]);

        Sum2[535]<=1^0^Co2[534];
        Co2[535]<=(1&0|(1|0)&Co2[534]);

        Sum2[536]<=1^0^Co2[535];
        Co2[536]<=(1&0|(1|0)&Co2[535]);

        Sum2[537]<=1^0^Co2[536];
        Co2[537]<=(1&0|(1|0)&Co2[536]);

        Sum2[538]<=1^0^Co2[537];
        Co2[538]<=(1&0|(1|0)&Co2[537]);

        Sum2[539]<=1^0^Co2[538];
        Co2[539]<=(1&0|(1|0)&Co2[538]);

        Sum2[540]<=1^0^Co2[539];
        Co2[540]<=(1&0|(1|0)&Co2[539]);

        Sum2[541]<=1^0^Co2[540];
        Co2[541]<=(1&0|(1|0)&Co2[540]);

        Sum2[542]<=1^0^Co2[541];
        Co2[542]<=(1&0|(1|0)&Co2[541]);

        Sum2[543]<=1^0^Co2[542];
        Co2[543]<=(1&0|(1|0)&Co2[542]);

        Sum2[544]<=1^0^Co2[543];
        Co2[544]<=(1&0|(1|0)&Co2[543]);

        Sum2[545]<=1^0^Co2[544];
        Co2[545]<=(1&0|(1|0)&Co2[544]);

        Sum2[546]<=1^0^Co2[545];
        Co2[546]<=(1&0|(1|0)&Co2[545]);

        Sum2[547]<=1^0^Co2[546];
        Co2[547]<=(1&0|(1|0)&Co2[546]);

        Sum2[548]<=1^0^Co2[547];
        Co2[548]<=(1&0|(1|0)&Co2[547]);

        Sum2[549]<=1^0^Co2[548];
        Co2[549]<=(1&0|(1|0)&Co2[548]);

        Sum2[550]<=1^0^Co2[549];
        Co2[550]<=(1&0|(1|0)&Co2[549]);

        Sum2[551]<=1^0^Co2[550];
        Co2[551]<=(1&0|(1|0)&Co2[550]);

        Sum2[552]<=1^0^Co2[551];
        Co2[552]<=(1&0|(1|0)&Co2[551]);

        Sum2[553]<=1^0^Co2[552];
        Co2[553]<=(1&0|(1|0)&Co2[552]);

        Sum2[554]<=1^0^Co2[553];
        Co2[554]<=(1&0|(1|0)&Co2[553]);

        Sum2[555]<=1^0^Co2[554];
        Co2[555]<=(1&0|(1|0)&Co2[554]);

        Sum2[556]<=1^0^Co2[555];
        Co2[556]<=(1&0|(1|0)&Co2[555]);

        Sum2[557]<=1^0^Co2[556];
        Co2[557]<=(1&0|(1|0)&Co2[556]);

        Sum2[558]<=1^0^Co2[557];
        Co2[558]<=(1&0|(1|0)&Co2[557]);

        Sum2[559]<=1^0^Co2[558];
        Co2[559]<=(1&0|(1|0)&Co2[558]);

        Sum2[560]<=1^0^Co2[559];
        Co2[560]<=(1&0|(1|0)&Co2[559]);

        Sum2[561]<=1^0^Co2[560];
        Co2[561]<=(1&0|(1|0)&Co2[560]);

        Sum2[562]<=1^0^Co2[561];
        Co2[562]<=(1&0|(1|0)&Co2[561]);

        Sum2[563]<=1^0^Co2[562];
        Co2[563]<=(1&0|(1|0)&Co2[562]);

        Sum2[564]<=1^0^Co2[563];
        Co2[564]<=(1&0|(1|0)&Co2[563]);

        Sum2[565]<=1^0^Co2[564];
        Co2[565]<=(1&0|(1|0)&Co2[564]);

        Sum2[566]<=1^0^Co2[565];
        Co2[566]<=(1&0|(1|0)&Co2[565]);

        Sum2[567]<=1^0^Co2[566];
        Co2[567]<=(1&0|(1|0)&Co2[566]);

        Sum2[568]<=1^0^Co2[567];
        Co2[568]<=(1&0|(1|0)&Co2[567]);

        Sum2[569]<=1^0^Co2[568];
        Co2[569]<=(1&0|(1|0)&Co2[568]);

        Sum2[570]<=1^0^Co2[569];
        Co2[570]<=(1&0|(1|0)&Co2[569]);

        Sum2[571]<=1^0^Co2[570];
        Co2[571]<=(1&0|(1|0)&Co2[570]);

        Sum2[572]<=1^0^Co2[571];
        Co2[572]<=(1&0|(1|0)&Co2[571]);

        Sum2[573]<=1^0^Co2[572];
        Co2[573]<=(1&0|(1|0)&Co2[572]);

        Sum2[574]<=1^0^Co2[573];
        Co2[574]<=(1&0|(1|0)&Co2[573]);

        Sum2[575]<=1^0^Co2[574];
        Co2[575]<=(1&0|(1|0)&Co2[574]);

        Sum2[576]<=1^0^Co2[575];
        Co2[576]<=(1&0|(1|0)&Co2[575]);

        Sum2[577]<=1^0^Co2[576];
        Co2[577]<=(1&0|(1|0)&Co2[576]);

        Sum2[578]<=1^0^Co2[577];
        Co2[578]<=(1&0|(1|0)&Co2[577]);

        Sum2[579]<=1^0^Co2[578];
        Co2[579]<=(1&0|(1|0)&Co2[578]);

        Sum2[580]<=1^0^Co2[579];
        Co2[580]<=(1&0|(1|0)&Co2[579]);

        Sum2[581]<=1^0^Co2[580];
        Co2[581]<=(1&0|(1|0)&Co2[580]);

        Sum2[582]<=1^0^Co2[581];
        Co2[582]<=(1&0|(1|0)&Co2[581]);

        Sum2[583]<=1^0^Co2[582];
        Co2[583]<=(1&0|(1|0)&Co2[582]);

        Sum2[584]<=1^0^Co2[583];
        Co2[584]<=(1&0|(1|0)&Co2[583]);

        Sum2[585]<=1^0^Co2[584];
        Co2[585]<=(1&0|(1|0)&Co2[584]);

        Sum2[586]<=1^0^Co2[585];
        Co2[586]<=(1&0|(1|0)&Co2[585]);

        Sum2[587]<=1^0^Co2[586];
        Co2[587]<=(1&0|(1|0)&Co2[586]);

        Sum2[588]<=1^0^Co2[587];
        Co2[588]<=(1&0|(1|0)&Co2[587]);

        Sum2[589]<=1^0^Co2[588];
        Co2[589]<=(1&0|(1|0)&Co2[588]);

        Sum2[590]<=1^0^Co2[589];
        Co2[590]<=(1&0|(1|0)&Co2[589]);

        Sum2[591]<=1^0^Co2[590];
        Co2[591]<=(1&0|(1|0)&Co2[590]);

        Sum2[592]<=1^0^Co2[591];
        Co2[592]<=(1&0|(1|0)&Co2[591]);

        Sum2[593]<=1^0^Co2[592];
        Co2[593]<=(1&0|(1|0)&Co2[592]);

        Sum2[594]<=1^0^Co2[593];
        Co2[594]<=(1&0|(1|0)&Co2[593]);

        Sum2[595]<=1^0^Co2[594];
        Co2[595]<=(1&0|(1|0)&Co2[594]);

        Sum2[596]<=1^0^Co2[595];
        Co2[596]<=(1&0|(1|0)&Co2[595]);

        Sum2[597]<=1^0^Co2[596];
        Co2[597]<=(1&0|(1|0)&Co2[596]);

        Sum2[598]<=1^0^Co2[597];
        Co2[598]<=(1&0|(1|0)&Co2[597]);

        Sum2[599]<=1^0^Co2[598];
        Co2[599]<=(1&0|(1|0)&Co2[598]);

        Sum2[600]<=1^0^Co2[599];
        Co2[600]<=(1&0|(1|0)&Co2[599]);

        Sum2[601]<=1^0^Co2[600];
        Co2[601]<=(1&0|(1|0)&Co2[600]);

        Sum2[602]<=1^0^Co2[601];
        Co2[602]<=(1&0|(1|0)&Co2[601]);

        Sum2[603]<=1^0^Co2[602];
        Co2[603]<=(1&0|(1|0)&Co2[602]);

        Sum2[604]<=1^0^Co2[603];
        Co2[604]<=(1&0|(1|0)&Co2[603]);

        Sum2[605]<=1^0^Co2[604];
        Co2[605]<=(1&0|(1|0)&Co2[604]);

        Sum2[606]<=1^0^Co2[605];
        Co2[606]<=(1&0|(1|0)&Co2[605]);

        Sum2[607]<=1^0^Co2[606];
        Co2[607]<=(1&0|(1|0)&Co2[606]);

        Sum2[608]<=1^0^Co2[607];
        Co2[608]<=(1&0|(1|0)&Co2[607]);

        Sum2[609]<=1^0^Co2[608];
        Co2[609]<=(1&0|(1|0)&Co2[608]);

        Sum2[610]<=1^0^Co2[609];
        Co2[610]<=(1&0|(1|0)&Co2[609]);

        Sum2[611]<=1^0^Co2[610];
        Co2[611]<=(1&0|(1|0)&Co2[610]);

        Sum2[612]<=1^0^Co2[611];
        Co2[612]<=(1&0|(1|0)&Co2[611]);

        Sum2[613]<=1^0^Co2[612];
        Co2[613]<=(1&0|(1|0)&Co2[612]);

        Sum2[614]<=1^0^Co2[613];
        Co2[614]<=(1&0|(1|0)&Co2[613]);

        Sum2[615]<=1^0^Co2[614];
        Co2[615]<=(1&0|(1|0)&Co2[614]);

        Sum2[616]<=1^0^Co2[615];
        Co2[616]<=(1&0|(1|0)&Co2[615]);

        Sum2[617]<=1^0^Co2[616];
        Co2[617]<=(1&0|(1|0)&Co2[616]);

        Sum2[618]<=1^0^Co2[617];
        Co2[618]<=(1&0|(1|0)&Co2[617]);

        Sum2[619]<=1^0^Co2[618];
        Co2[619]<=(1&0|(1|0)&Co2[618]);

        Sum2[620]<=1^0^Co2[619];
        Co2[620]<=(1&0|(1|0)&Co2[619]);

        Sum2[621]<=1^0^Co2[620];
        Co2[621]<=(1&0|(1|0)&Co2[620]);

        Sum2[622]<=1^0^Co2[621];
        Co2[622]<=(1&0|(1|0)&Co2[621]);

        Sum2[623]<=1^0^Co2[622];
        Co2[623]<=(1&0|(1|0)&Co2[622]);

        Sum2[624]<=1^0^Co2[623];
        Co2[624]<=(1&0|(1|0)&Co2[623]);

        Sum2[625]<=1^0^Co2[624];
        Co2[625]<=(1&0|(1|0)&Co2[624]);

        Sum2[626]<=1^0^Co2[625];
        Co2[626]<=(1&0|(1|0)&Co2[625]);

        Sum2[627]<=1^0^Co2[626];
        Co2[627]<=(1&0|(1|0)&Co2[626]);

        Sum2[628]<=1^0^Co2[627];
        Co2[628]<=(1&0|(1|0)&Co2[627]);

        Sum2[629]<=1^0^Co2[628];
        Co2[629]<=(1&0|(1|0)&Co2[628]);

        Sum2[630]<=1^0^Co2[629];
        Co2[630]<=(1&0|(1|0)&Co2[629]);

        Sum2[631]<=1^0^Co2[630];
        Co2[631]<=(1&0|(1|0)&Co2[630]);

        Sum2[632]<=1^0^Co2[631];
        Co2[632]<=(1&0|(1|0)&Co2[631]);

        Sum2[633]<=1^0^Co2[632];
        Co2[633]<=(1&0|(1|0)&Co2[632]);

        Sum2[634]<=1^0^Co2[633];
        Co2[634]<=(1&0|(1|0)&Co2[633]);

        Sum2[635]<=1^0^Co2[634];
        Co2[635]<=(1&0|(1|0)&Co2[634]);

        Sum2[636]<=1^0^Co2[635];
        Co2[636]<=(1&0|(1|0)&Co2[635]);

        Sum2[637]<=1^0^Co2[636];
        Co2[637]<=(1&0|(1|0)&Co2[636]);

        Sum2[638]<=1^0^Co2[637];
        Co2[638]<=(1&0|(1|0)&Co2[637]);

        Sum2[639]<=1^0^Co2[638];
        Co2[639]<=(1&0|(1|0)&Co2[638]);

        Sum2[640]<=1^0^Co2[639];
        Co2[640]<=(1&0|(1|0)&Co2[639]);

        Sum2[641]<=1^0^Co2[640];
        Co2[641]<=(1&0|(1|0)&Co2[640]);

        Sum2[642]<=1^0^Co2[641];
        Co2[642]<=(1&0|(1|0)&Co2[641]);

        Sum2[643]<=1^0^Co2[642];
        Co2[643]<=(1&0|(1|0)&Co2[642]);

        Sum2[644]<=1^0^Co2[643];
        Co2[644]<=(1&0|(1|0)&Co2[643]);

        Sum2[645]<=1^0^Co2[644];
        Co2[645]<=(1&0|(1|0)&Co2[644]);

        Sum2[646]<=1^0^Co2[645];
        Co2[646]<=(1&0|(1|0)&Co2[645]);

        Sum2[647]<=1^0^Co2[646];
        Co2[647]<=(1&0|(1|0)&Co2[646]);

        Sum2[648]<=1^0^Co2[647];
        Co2[648]<=(1&0|(1|0)&Co2[647]);

        Sum2[649]<=1^0^Co2[648];
        Co2[649]<=(1&0|(1|0)&Co2[648]);

        Sum2[650]<=1^0^Co2[649];
        Co2[650]<=(1&0|(1|0)&Co2[649]);

        Sum2[651]<=1^0^Co2[650];
        Co2[651]<=(1&0|(1|0)&Co2[650]);

        Sum2[652]<=1^0^Co2[651];
        Co2[652]<=(1&0|(1|0)&Co2[651]);

        Sum2[653]<=1^0^Co2[652];
        Co2[653]<=(1&0|(1|0)&Co2[652]);

        Sum2[654]<=1^0^Co2[653];
        Co2[654]<=(1&0|(1|0)&Co2[653]);

        Sum2[655]<=1^0^Co2[654];
        Co2[655]<=(1&0|(1|0)&Co2[654]);

        Sum2[656]<=1^0^Co2[655];
        Co2[656]<=(1&0|(1|0)&Co2[655]);

        Sum2[657]<=1^0^Co2[656];
        Co2[657]<=(1&0|(1|0)&Co2[656]);

        Sum2[658]<=1^0^Co2[657];
        Co2[658]<=(1&0|(1|0)&Co2[657]);

        Sum2[659]<=1^0^Co2[658];
        Co2[659]<=(1&0|(1|0)&Co2[658]);

        Sum2[660]<=1^0^Co2[659];
        Co2[660]<=(1&0|(1|0)&Co2[659]);

        Sum2[661]<=1^0^Co2[660];
        Co2[661]<=(1&0|(1|0)&Co2[660]);

        Sum2[662]<=1^0^Co2[661];
        Co2[662]<=(1&0|(1|0)&Co2[661]);

        Sum2[663]<=1^0^Co2[662];
        Co2[663]<=(1&0|(1|0)&Co2[662]);

        Sum2[664]<=1^0^Co2[663];
        Co2[664]<=(1&0|(1|0)&Co2[663]);

        Sum2[665]<=1^0^Co2[664];
        Co2[665]<=(1&0|(1|0)&Co2[664]);

        Sum2[666]<=1^0^Co2[665];
        Co2[666]<=(1&0|(1|0)&Co2[665]);

        Sum2[667]<=1^0^Co2[666];
        Co2[667]<=(1&0|(1|0)&Co2[666]);

        Sum2[668]<=1^0^Co2[667];
        Co2[668]<=(1&0|(1|0)&Co2[667]);

        Sum2[669]<=1^0^Co2[668];
        Co2[669]<=(1&0|(1|0)&Co2[668]);

        Sum2[670]<=1^0^Co2[669];
        Co2[670]<=(1&0|(1|0)&Co2[669]);

        Sum2[671]<=1^0^Co2[670];
        Co2[671]<=(1&0|(1|0)&Co2[670]);

        Sum2[672]<=1^0^Co2[671];
        Co2[672]<=(1&0|(1|0)&Co2[671]);

        Sum2[673]<=1^0^Co2[672];
        Co2[673]<=(1&0|(1|0)&Co2[672]);

        Sum2[674]<=1^0^Co2[673];
        Co2[674]<=(1&0|(1|0)&Co2[673]);

        Sum2[675]<=1^0^Co2[674];
        Co2[675]<=(1&0|(1|0)&Co2[674]);

        Sum2[676]<=1^0^Co2[675];
        Co2[676]<=(1&0|(1|0)&Co2[675]);

        Sum2[677]<=1^0^Co2[676];
        Co2[677]<=(1&0|(1|0)&Co2[676]);

        Sum2[678]<=1^0^Co2[677];
        Co2[678]<=(1&0|(1|0)&Co2[677]);

        Sum2[679]<=1^0^Co2[678];
        Co2[679]<=(1&0|(1|0)&Co2[678]);

        Sum2[680]<=1^0^Co2[679];
        Co2[680]<=(1&0|(1|0)&Co2[679]);

        Sum2[681]<=1^0^Co2[680];
        Co2[681]<=(1&0|(1|0)&Co2[680]);

        Sum2[682]<=1^0^Co2[681];
        Co2[682]<=(1&0|(1|0)&Co2[681]);

        Sum2[683]<=1^0^Co2[682];
        Co2[683]<=(1&0|(1|0)&Co2[682]);

        Sum2[684]<=1^0^Co2[683];
        Co2[684]<=(1&0|(1|0)&Co2[683]);

        Sum2[685]<=1^0^Co2[684];
        Co2[685]<=(1&0|(1|0)&Co2[684]);

        Sum2[686]<=1^0^Co2[685];
        Co2[686]<=(1&0|(1|0)&Co2[685]);

        Sum2[687]<=1^0^Co2[686];
        Co2[687]<=(1&0|(1|0)&Co2[686]);

        Sum2[688]<=1^0^Co2[687];
        Co2[688]<=(1&0|(1|0)&Co2[687]);

        Sum2[689]<=1^0^Co2[688];
        Co2[689]<=(1&0|(1|0)&Co2[688]);

        Sum2[690]<=1^0^Co2[689];
        Co2[690]<=(1&0|(1|0)&Co2[689]);

        Sum2[691]<=1^0^Co2[690];
        Co2[691]<=(1&0|(1|0)&Co2[690]);

        Sum2[692]<=1^0^Co2[691];
        Co2[692]<=(1&0|(1|0)&Co2[691]);

        Sum2[693]<=1^0^Co2[692];
        Co2[693]<=(1&0|(1|0)&Co2[692]);

        Sum2[694]<=1^0^Co2[693];
        Co2[694]<=(1&0|(1|0)&Co2[693]);

        Sum2[695]<=1^0^Co2[694];
        Co2[695]<=(1&0|(1|0)&Co2[694]);

        Sum2[696]<=1^0^Co2[695];
        Co2[696]<=(1&0|(1|0)&Co2[695]);

        Sum2[697]<=1^0^Co2[696];
        Co2[697]<=(1&0|(1|0)&Co2[696]);

        Sum2[698]<=1^0^Co2[697];
        Co2[698]<=(1&0|(1|0)&Co2[697]);

        Sum2[699]<=1^0^Co2[698];
        Co2[699]<=(1&0|(1|0)&Co2[698]);

        Sum2[700]<=1^0^Co2[699];
        Co2[700]<=(1&0|(1|0)&Co2[699]);

        Sum2[701]<=1^0^Co2[700];
        Co2[701]<=(1&0|(1|0)&Co2[700]);

        Sum2[702]<=1^0^Co2[701];
        Co2[702]<=(1&0|(1|0)&Co2[701]);

        Sum2[703]<=1^0^Co2[702];
        Co2[703]<=(1&0|(1|0)&Co2[702]);

        Sum2[704]<=1^0^Co2[703];
        Co2[704]<=(1&0|(1|0)&Co2[703]);

        Sum2[705]<=1^0^Co2[704];
        Co2[705]<=(1&0|(1|0)&Co2[704]);

        Sum2[706]<=1^0^Co2[705];
        Co2[706]<=(1&0|(1|0)&Co2[705]);

        Sum2[707]<=1^0^Co2[706];
        Co2[707]<=(1&0|(1|0)&Co2[706]);

        Sum2[708]<=1^0^Co2[707];
        Co2[708]<=(1&0|(1|0)&Co2[707]);

        Sum2[709]<=1^0^Co2[708];
        Co2[709]<=(1&0|(1|0)&Co2[708]);

        Sum2[710]<=1^0^Co2[709];
        Co2[710]<=(1&0|(1|0)&Co2[709]);

        Sum2[711]<=1^0^Co2[710];
        Co2[711]<=(1&0|(1|0)&Co2[710]);

        Sum2[712]<=1^0^Co2[711];
        Co2[712]<=(1&0|(1|0)&Co2[711]);

        Sum2[713]<=1^0^Co2[712];
        Co2[713]<=(1&0|(1|0)&Co2[712]);

        Sum2[714]<=1^0^Co2[713];
        Co2[714]<=(1&0|(1|0)&Co2[713]);

        Sum2[715]<=1^0^Co2[714];
        Co2[715]<=(1&0|(1|0)&Co2[714]);

        Sum2[716]<=1^0^Co2[715];
        Co2[716]<=(1&0|(1|0)&Co2[715]);

        Sum2[717]<=1^0^Co2[716];
        Co2[717]<=(1&0|(1|0)&Co2[716]);

        Sum2[718]<=1^0^Co2[717];
        Co2[718]<=(1&0|(1|0)&Co2[717]);

        Sum2[719]<=1^0^Co2[718];
        Co2[719]<=(1&0|(1|0)&Co2[718]);

        Sum2[720]<=1^0^Co2[719];
        Co2[720]<=(1&0|(1|0)&Co2[719]);

        Sum2[721]<=1^0^Co2[720];
        Co2[721]<=(1&0|(1|0)&Co2[720]);

        Sum2[722]<=1^0^Co2[721];
        Co2[722]<=(1&0|(1|0)&Co2[721]);

        Sum2[723]<=1^0^Co2[722];
        Co2[723]<=(1&0|(1|0)&Co2[722]);

        Sum2[724]<=1^0^Co2[723];
        Co2[724]<=(1&0|(1|0)&Co2[723]);

        Sum2[725]<=1^0^Co2[724];
        Co2[725]<=(1&0|(1|0)&Co2[724]);

        Sum2[726]<=1^0^Co2[725];
        Co2[726]<=(1&0|(1|0)&Co2[725]);

        Sum2[727]<=1^0^Co2[726];
        Co2[727]<=(1&0|(1|0)&Co2[726]);

        Sum2[728]<=1^0^Co2[727];
        Co2[728]<=(1&0|(1|0)&Co2[727]);

        Sum2[729]<=1^0^Co2[728];
        Co2[729]<=(1&0|(1|0)&Co2[728]);

        Sum2[730]<=1^0^Co2[729];
        Co2[730]<=(1&0|(1|0)&Co2[729]);

        Sum2[731]<=1^0^Co2[730];
        Co2[731]<=(1&0|(1|0)&Co2[730]);

        Sum2[732]<=1^0^Co2[731];
        Co2[732]<=(1&0|(1|0)&Co2[731]);

        Sum2[733]<=1^0^Co2[732];
        Co2[733]<=(1&0|(1|0)&Co2[732]);

        Sum2[734]<=1^0^Co2[733];
        Co2[734]<=(1&0|(1|0)&Co2[733]);

        Sum2[735]<=1^0^Co2[734];
        Co2[735]<=(1&0|(1|0)&Co2[734]);

        Sum2[736]<=1^0^Co2[735];
        Co2[736]<=(1&0|(1|0)&Co2[735]);

        Sum2[737]<=1^0^Co2[736];
        Co2[737]<=(1&0|(1|0)&Co2[736]);

        Sum2[738]<=1^0^Co2[737];
        Co2[738]<=(1&0|(1|0)&Co2[737]);

        Sum2[739]<=1^0^Co2[738];
        Co2[739]<=(1&0|(1|0)&Co2[738]);

        Sum2[740]<=1^0^Co2[739];
        Co2[740]<=(1&0|(1|0)&Co2[739]);

        Sum2[741]<=1^0^Co2[740];
        Co2[741]<=(1&0|(1|0)&Co2[740]);

        Sum2[742]<=1^0^Co2[741];
        Co2[742]<=(1&0|(1|0)&Co2[741]);

        Sum2[743]<=1^0^Co2[742];
        Co2[743]<=(1&0|(1|0)&Co2[742]);

        Sum2[744]<=1^0^Co2[743];
        Co2[744]<=(1&0|(1|0)&Co2[743]);

        Sum2[745]<=1^0^Co2[744];
        Co2[745]<=(1&0|(1|0)&Co2[744]);

        Sum2[746]<=1^0^Co2[745];
        Co2[746]<=(1&0|(1|0)&Co2[745]);

        Sum2[747]<=1^0^Co2[746];
        Co2[747]<=(1&0|(1|0)&Co2[746]);

        Sum2[748]<=1^0^Co2[747];
        Co2[748]<=(1&0|(1|0)&Co2[747]);

        Sum2[749]<=1^0^Co2[748];
        Co2[749]<=(1&0|(1|0)&Co2[748]);

        Sum2[750]<=1^0^Co2[749];
        Co2[750]<=(1&0|(1|0)&Co2[749]);

        Sum2[751]<=1^0^Co2[750];
        Co2[751]<=(1&0|(1|0)&Co2[750]);

        Sum2[752]<=1^0^Co2[751];
        Co2[752]<=(1&0|(1|0)&Co2[751]);

        Sum2[753]<=1^0^Co2[752];
        Co2[753]<=(1&0|(1|0)&Co2[752]);

        Sum2[754]<=1^0^Co2[753];
        Co2[754]<=(1&0|(1|0)&Co2[753]);

        Sum2[755]<=1^0^Co2[754];
        Co2[755]<=(1&0|(1|0)&Co2[754]);

        Sum2[756]<=1^0^Co2[755];
        Co2[756]<=(1&0|(1|0)&Co2[755]);

        Sum2[757]<=1^0^Co2[756];
        Co2[757]<=(1&0|(1|0)&Co2[756]);

        Sum2[758]<=1^0^Co2[757];
        Co2[758]<=(1&0|(1|0)&Co2[757]);

        Sum2[759]<=1^0^Co2[758];
        Co2[759]<=(1&0|(1|0)&Co2[758]);

        Sum2[760]<=1^0^Co2[759];
        Co2[760]<=(1&0|(1|0)&Co2[759]);

        Sum2[761]<=1^0^Co2[760];
        Co2[761]<=(1&0|(1|0)&Co2[760]);

        Sum2[762]<=1^0^Co2[761];
        Co2[762]<=(1&0|(1|0)&Co2[761]);

        Sum2[763]<=1^0^Co2[762];
        Co2[763]<=(1&0|(1|0)&Co2[762]);

        Sum2[764]<=1^0^Co2[763];
        Co2[764]<=(1&0|(1|0)&Co2[763]);

        Sum2[765]<=1^0^Co2[764];
        Co2[765]<=(1&0|(1|0)&Co2[764]);

        Sum2[766]<=1^0^Co2[765];
        Co2[766]<=(1&0|(1|0)&Co2[765]);

        Sum2[767]<=1^0^Co2[766];
        Co2[767]<=(1&0|(1|0)&Co2[766]);

        Sum2[768]<=1^0^Co2[767];
        Co2[768]<=(1&0|(1|0)&Co2[767]);

        Sum2[769]<=1^0^Co2[768];
        Co2[769]<=(1&0|(1|0)&Co2[768]);

        Sum2[770]<=1^0^Co2[769];
        Co2[770]<=(1&0|(1|0)&Co2[769]);

        Sum2[771]<=1^0^Co2[770];
        Co2[771]<=(1&0|(1|0)&Co2[770]);

        Sum2[772]<=1^0^Co2[771];
        Co2[772]<=(1&0|(1|0)&Co2[771]);

        Sum2[773]<=1^0^Co2[772];
        Co2[773]<=(1&0|(1|0)&Co2[772]);

        Sum2[774]<=1^0^Co2[773];
        Co2[774]<=(1&0|(1|0)&Co2[773]);

        Sum2[775]<=1^0^Co2[774];
        Co2[775]<=(1&0|(1|0)&Co2[774]);

        Sum2[776]<=1^0^Co2[775];
        Co2[776]<=(1&0|(1|0)&Co2[775]);

        Sum2[777]<=1^0^Co2[776];
        Co2[777]<=(1&0|(1|0)&Co2[776]);

        Sum2[778]<=1^0^Co2[777];
        Co2[778]<=(1&0|(1|0)&Co2[777]);

        Sum2[779]<=1^0^Co2[778];
        Co2[779]<=(1&0|(1|0)&Co2[778]);

        Sum2[780]<=1^0^Co2[779];
        Co2[780]<=(1&0|(1|0)&Co2[779]);

        Sum2[781]<=1^0^Co2[780];
        Co2[781]<=(1&0|(1|0)&Co2[780]);

        Sum2[782]<=1^0^Co2[781];
        Co2[782]<=(1&0|(1|0)&Co2[781]);

        Sum2[783]<=1^0^Co2[782];
        Co2[783]<=(1&0|(1|0)&Co2[782]);

        Sum2[784]<=1^0^Co2[783];
        Co2[784]<=(1&0|(1|0)&Co2[783]);

        Sum2[785]<=1^0^Co2[784];
        Co2[785]<=(1&0|(1|0)&Co2[784]);

        Sum2[786]<=1^0^Co2[785];
        Co2[786]<=(1&0|(1|0)&Co2[785]);

        Sum2[787]<=1^0^Co2[786];
        Co2[787]<=(1&0|(1|0)&Co2[786]);

        Sum2[788]<=1^0^Co2[787];
        Co2[788]<=(1&0|(1|0)&Co2[787]);

        Sum2[789]<=1^0^Co2[788];
        Co2[789]<=(1&0|(1|0)&Co2[788]);

        Sum2[790]<=1^0^Co2[789];
        Co2[790]<=(1&0|(1|0)&Co2[789]);

        Sum2[791]<=1^0^Co2[790];
        Co2[791]<=(1&0|(1|0)&Co2[790]);

        Sum2[792]<=1^0^Co2[791];
        Co2[792]<=(1&0|(1|0)&Co2[791]);

        Sum2[793]<=1^0^Co2[792];
        Co2[793]<=(1&0|(1|0)&Co2[792]);

        Sum2[794]<=1^0^Co2[793];
        Co2[794]<=(1&0|(1|0)&Co2[793]);

        Sum2[795]<=1^0^Co2[794];
        Co2[795]<=(1&0|(1|0)&Co2[794]);

        Sum2[796]<=1^0^Co2[795];
        Co2[796]<=(1&0|(1|0)&Co2[795]);

        Sum2[797]<=1^0^Co2[796];
        Co2[797]<=(1&0|(1|0)&Co2[796]);

        Sum2[798]<=1^0^Co2[797];
        Co2[798]<=(1&0|(1|0)&Co2[797]);

        Sum2[799]<=1^0^Co2[798];
        Co2[799]<=(1&0|(1|0)&Co2[798]);

        Sum2[800]<=1^0^Co2[799];
        Co2[800]<=(1&0|(1|0)&Co2[799]);

        Sum2[801]<=1^0^Co2[800];
        Co2[801]<=(1&0|(1|0)&Co2[800]);

        Sum2[802]<=1^0^Co2[801];
        Co2[802]<=(1&0|(1|0)&Co2[801]);

        Sum2[803]<=1^0^Co2[802];
        Co2[803]<=(1&0|(1|0)&Co2[802]);

        Sum2[804]<=1^0^Co2[803];
        Co2[804]<=(1&0|(1|0)&Co2[803]);

        Sum2[805]<=1^0^Co2[804];
        Co2[805]<=(1&0|(1|0)&Co2[804]);

        Sum2[806]<=1^0^Co2[805];
        Co2[806]<=(1&0|(1|0)&Co2[805]);

        Sum2[807]<=1^0^Co2[806];
        Co2[807]<=(1&0|(1|0)&Co2[806]);

        Sum2[808]<=1^0^Co2[807];
        Co2[808]<=(1&0|(1|0)&Co2[807]);

        Sum2[809]<=1^0^Co2[808];
        Co2[809]<=(1&0|(1|0)&Co2[808]);

        Sum2[810]<=1^0^Co2[809];
        Co2[810]<=(1&0|(1|0)&Co2[809]);

        Sum2[811]<=1^0^Co2[810];
        Co2[811]<=(1&0|(1|0)&Co2[810]);

        Sum2[812]<=1^0^Co2[811];
        Co2[812]<=(1&0|(1|0)&Co2[811]);

        Sum2[813]<=1^0^Co2[812];
        Co2[813]<=(1&0|(1|0)&Co2[812]);

        Sum2[814]<=1^0^Co2[813];
        Co2[814]<=(1&0|(1|0)&Co2[813]);

        Sum2[815]<=1^0^Co2[814];
        Co2[815]<=(1&0|(1|0)&Co2[814]);

        Sum2[816]<=1^0^Co2[815];
        Co2[816]<=(1&0|(1|0)&Co2[815]);

        Sum2[817]<=1^0^Co2[816];
        Co2[817]<=(1&0|(1|0)&Co2[816]);

        Sum2[818]<=1^0^Co2[817];
        Co2[818]<=(1&0|(1|0)&Co2[817]);

        Sum2[819]<=1^0^Co2[818];
        Co2[819]<=(1&0|(1|0)&Co2[818]);

        Sum2[820]<=1^0^Co2[819];
        Co2[820]<=(1&0|(1|0)&Co2[819]);

        Sum2[821]<=1^0^Co2[820];
        Co2[821]<=(1&0|(1|0)&Co2[820]);

        Sum2[822]<=1^0^Co2[821];
        Co2[822]<=(1&0|(1|0)&Co2[821]);

        Sum2[823]<=1^0^Co2[822];
        Co2[823]<=(1&0|(1|0)&Co2[822]);

        Sum2[824]<=1^0^Co2[823];
        Co2[824]<=(1&0|(1|0)&Co2[823]);

        Sum2[825]<=1^0^Co2[824];
        Co2[825]<=(1&0|(1|0)&Co2[824]);

        Sum2[826]<=1^0^Co2[825];
        Co2[826]<=(1&0|(1|0)&Co2[825]);

        Sum2[827]<=1^0^Co2[826];
        Co2[827]<=(1&0|(1|0)&Co2[826]);

        Sum2[828]<=1^0^Co2[827];
        Co2[828]<=(1&0|(1|0)&Co2[827]);

        Sum2[829]<=1^0^Co2[828];
        Co2[829]<=(1&0|(1|0)&Co2[828]);

        Sum2[830]<=1^0^Co2[829];
        Co2[830]<=(1&0|(1|0)&Co2[829]);

        Sum2[831]<=1^0^Co2[830];
        Co2[831]<=(1&0|(1|0)&Co2[830]);

        Sum2[832]<=1^0^Co2[831];
        Co2[832]<=(1&0|(1|0)&Co2[831]);

        Sum2[833]<=1^0^Co2[832];
        Co2[833]<=(1&0|(1|0)&Co2[832]);

        Sum2[834]<=1^0^Co2[833];
        Co2[834]<=(1&0|(1|0)&Co2[833]);

        Sum2[835]<=1^0^Co2[834];
        Co2[835]<=(1&0|(1|0)&Co2[834]);

        Sum2[836]<=1^0^Co2[835];
        Co2[836]<=(1&0|(1|0)&Co2[835]);

        Sum2[837]<=1^0^Co2[836];
        Co2[837]<=(1&0|(1|0)&Co2[836]);

        Sum2[838]<=1^0^Co2[837];
        Co2[838]<=(1&0|(1|0)&Co2[837]);

        Sum2[839]<=1^0^Co2[838];
        Co2[839]<=(1&0|(1|0)&Co2[838]);

        Sum2[840]<=1^0^Co2[839];
        Co2[840]<=(1&0|(1|0)&Co2[839]);

        Sum2[841]<=1^0^Co2[840];
        Co2[841]<=(1&0|(1|0)&Co2[840]);

        Sum2[842]<=1^0^Co2[841];
        Co2[842]<=(1&0|(1|0)&Co2[841]);

        Sum2[843]<=1^0^Co2[842];
        Co2[843]<=(1&0|(1|0)&Co2[842]);

        Sum2[844]<=1^0^Co2[843];
        Co2[844]<=(1&0|(1|0)&Co2[843]);

        Sum2[845]<=1^0^Co2[844];
        Co2[845]<=(1&0|(1|0)&Co2[844]);

        Sum2[846]<=1^0^Co2[845];
        Co2[846]<=(1&0|(1|0)&Co2[845]);

        Sum2[847]<=1^0^Co2[846];
        Co2[847]<=(1&0|(1|0)&Co2[846]);

        Sum2[848]<=1^0^Co2[847];
        Co2[848]<=(1&0|(1|0)&Co2[847]);

        Sum2[849]<=1^0^Co2[848];
        Co2[849]<=(1&0|(1|0)&Co2[848]);

        Sum2[850]<=1^0^Co2[849];
        Co2[850]<=(1&0|(1|0)&Co2[849]);

        Sum2[851]<=1^0^Co2[850];
        Co2[851]<=(1&0|(1|0)&Co2[850]);

        Sum2[852]<=1^0^Co2[851];
        Co2[852]<=(1&0|(1|0)&Co2[851]);

        Sum2[853]<=1^0^Co2[852];
        Co2[853]<=(1&0|(1|0)&Co2[852]);

        Sum2[854]<=1^0^Co2[853];
        Co2[854]<=(1&0|(1|0)&Co2[853]);

        Sum2[855]<=1^0^Co2[854];
        Co2[855]<=(1&0|(1|0)&Co2[854]);

        Sum2[856]<=1^0^Co2[855];
        Co2[856]<=(1&0|(1|0)&Co2[855]);

        Sum2[857]<=1^0^Co2[856];
        Co2[857]<=(1&0|(1|0)&Co2[856]);

        Sum2[858]<=1^0^Co2[857];
        Co2[858]<=(1&0|(1|0)&Co2[857]);

        Sum2[859]<=1^0^Co2[858];
        Co2[859]<=(1&0|(1|0)&Co2[858]);

        Sum2[860]<=1^0^Co2[859];
        Co2[860]<=(1&0|(1|0)&Co2[859]);

        Sum2[861]<=1^0^Co2[860];
        Co2[861]<=(1&0|(1|0)&Co2[860]);

        Sum2[862]<=1^0^Co2[861];
        Co2[862]<=(1&0|(1|0)&Co2[861]);

        Sum2[863]<=1^0^Co2[862];
        Co2[863]<=(1&0|(1|0)&Co2[862]);

        Sum2[864]<=1^0^Co2[863];
        Co2[864]<=(1&0|(1|0)&Co2[863]);

        Sum2[865]<=1^0^Co2[864];
        Co2[865]<=(1&0|(1|0)&Co2[864]);

        Sum2[866]<=1^0^Co2[865];
        Co2[866]<=(1&0|(1|0)&Co2[865]);

        Sum2[867]<=1^0^Co2[866];
        Co2[867]<=(1&0|(1|0)&Co2[866]);

        Sum2[868]<=1^0^Co2[867];
        Co2[868]<=(1&0|(1|0)&Co2[867]);

        Sum2[869]<=1^0^Co2[868];
        Co2[869]<=(1&0|(1|0)&Co2[868]);

        Sum2[870]<=1^0^Co2[869];
        Co2[870]<=(1&0|(1|0)&Co2[869]);

        Sum2[871]<=1^0^Co2[870];
        Co2[871]<=(1&0|(1|0)&Co2[870]);

        Sum2[872]<=1^0^Co2[871];
        Co2[872]<=(1&0|(1|0)&Co2[871]);

        Sum2[873]<=1^0^Co2[872];
        Co2[873]<=(1&0|(1|0)&Co2[872]);

        Sum2[874]<=1^0^Co2[873];
        Co2[874]<=(1&0|(1|0)&Co2[873]);

        Sum2[875]<=1^0^Co2[874];
        Co2[875]<=(1&0|(1|0)&Co2[874]);

        Sum2[876]<=1^0^Co2[875];
        Co2[876]<=(1&0|(1|0)&Co2[875]);

        Sum2[877]<=1^0^Co2[876];
        Co2[877]<=(1&0|(1|0)&Co2[876]);

        Sum2[878]<=1^0^Co2[877];
        Co2[878]<=(1&0|(1|0)&Co2[877]);

        Sum2[879]<=1^0^Co2[878];
        Co2[879]<=(1&0|(1|0)&Co2[878]);

        Sum2[880]<=1^0^Co2[879];
        Co2[880]<=(1&0|(1|0)&Co2[879]);

        Sum2[881]<=1^0^Co2[880];
        Co2[881]<=(1&0|(1|0)&Co2[880]);

        Sum2[882]<=1^0^Co2[881];
        Co2[882]<=(1&0|(1|0)&Co2[881]);

        Sum2[883]<=1^0^Co2[882];
        Co2[883]<=(1&0|(1|0)&Co2[882]);

        Sum2[884]<=1^0^Co2[883];
        Co2[884]<=(1&0|(1|0)&Co2[883]);

        Sum2[885]<=1^0^Co2[884];
        Co2[885]<=(1&0|(1|0)&Co2[884]);

        Sum2[886]<=1^0^Co2[885];
        Co2[886]<=(1&0|(1|0)&Co2[885]);

        Sum2[887]<=1^0^Co2[886];
        Co2[887]<=(1&0|(1|0)&Co2[886]);

        Sum2[888]<=1^0^Co2[887];
        Co2[888]<=(1&0|(1|0)&Co2[887]);

        Sum2[889]<=1^0^Co2[888];
        Co2[889]<=(1&0|(1|0)&Co2[888]);

        Sum2[890]<=1^0^Co2[889];
        Co2[890]<=(1&0|(1|0)&Co2[889]);

        Sum2[891]<=1^0^Co2[890];
        Co2[891]<=(1&0|(1|0)&Co2[890]);

        Sum2[892]<=1^0^Co2[891];
        Co2[892]<=(1&0|(1|0)&Co2[891]);

        Sum2[893]<=1^0^Co2[892];
        Co2[893]<=(1&0|(1|0)&Co2[892]);

        Sum2[894]<=1^0^Co2[893];
        Co2[894]<=(1&0|(1|0)&Co2[893]);

        Sum2[895]<=1^0^Co2[894];
        Co2[895]<=(1&0|(1|0)&Co2[894]);

        Sum2[896]<=1^0^Co2[895];
        Co2[896]<=(1&0|(1|0)&Co2[895]);

        Sum2[897]<=1^0^Co2[896];
        Co2[897]<=(1&0|(1|0)&Co2[896]);

        Sum2[898]<=1^0^Co2[897];
        Co2[898]<=(1&0|(1|0)&Co2[897]);

        Sum2[899]<=1^0^Co2[898];
        Co2[899]<=(1&0|(1|0)&Co2[898]);

        Sum2[900]<=1^0^Co2[899];
        Co2[900]<=(1&0|(1|0)&Co2[899]);

        Sum2[901]<=1^0^Co2[900];
        Co2[901]<=(1&0|(1|0)&Co2[900]);

        Sum2[902]<=1^0^Co2[901];
        Co2[902]<=(1&0|(1|0)&Co2[901]);

        Sum2[903]<=1^0^Co2[902];
        Co2[903]<=(1&0|(1|0)&Co2[902]);

        Sum2[904]<=1^0^Co2[903];
        Co2[904]<=(1&0|(1|0)&Co2[903]);

        Sum2[905]<=1^0^Co2[904];
        Co2[905]<=(1&0|(1|0)&Co2[904]);

        Sum2[906]<=1^0^Co2[905];
        Co2[906]<=(1&0|(1|0)&Co2[905]);

        Sum2[907]<=1^0^Co2[906];
        Co2[907]<=(1&0|(1|0)&Co2[906]);

        Sum2[908]<=1^0^Co2[907];
        Co2[908]<=(1&0|(1|0)&Co2[907]);

        Sum2[909]<=1^0^Co2[908];
        Co2[909]<=(1&0|(1|0)&Co2[908]);

        Sum2[910]<=1^0^Co2[909];
        Co2[910]<=(1&0|(1|0)&Co2[909]);

        Sum2[911]<=1^0^Co2[910];
        Co2[911]<=(1&0|(1|0)&Co2[910]);

        Sum2[912]<=1^0^Co2[911];
        Co2[912]<=(1&0|(1|0)&Co2[911]);

        Sum2[913]<=1^0^Co2[912];
        Co2[913]<=(1&0|(1|0)&Co2[912]);

        Sum2[914]<=1^0^Co2[913];
        Co2[914]<=(1&0|(1|0)&Co2[913]);

        Sum2[915]<=1^0^Co2[914];
        Co2[915]<=(1&0|(1|0)&Co2[914]);

        Sum2[916]<=1^0^Co2[915];
        Co2[916]<=(1&0|(1|0)&Co2[915]);

        Sum2[917]<=1^0^Co2[916];
        Co2[917]<=(1&0|(1|0)&Co2[916]);

        Sum2[918]<=1^0^Co2[917];
        Co2[918]<=(1&0|(1|0)&Co2[917]);

        Sum2[919]<=1^0^Co2[918];
        Co2[919]<=(1&0|(1|0)&Co2[918]);

        Sum2[920]<=1^0^Co2[919];
        Co2[920]<=(1&0|(1|0)&Co2[919]);

        Sum2[921]<=1^0^Co2[920];
        Co2[921]<=(1&0|(1|0)&Co2[920]);

        Sum2[922]<=1^0^Co2[921];
        Co2[922]<=(1&0|(1|0)&Co2[921]);

        Sum2[923]<=1^0^Co2[922];
        Co2[923]<=(1&0|(1|0)&Co2[922]);

        Sum2[924]<=1^0^Co2[923];
        Co2[924]<=(1&0|(1|0)&Co2[923]);

        Sum2[925]<=1^0^Co2[924];
        Co2[925]<=(1&0|(1|0)&Co2[924]);

        Sum2[926]<=1^0^Co2[925];
        Co2[926]<=(1&0|(1|0)&Co2[925]);

        Sum2[927]<=1^0^Co2[926];
        Co2[927]<=(1&0|(1|0)&Co2[926]);

        Sum2[928]<=1^0^Co2[927];
        Co2[928]<=(1&0|(1|0)&Co2[927]);

        Sum2[929]<=1^0^Co2[928];
        Co2[929]<=(1&0|(1|0)&Co2[928]);

        Sum2[930]<=1^0^Co2[929];
        Co2[930]<=(1&0|(1|0)&Co2[929]);

        Sum2[931]<=1^0^Co2[930];
        Co2[931]<=(1&0|(1|0)&Co2[930]);

        Sum2[932]<=1^0^Co2[931];
        Co2[932]<=(1&0|(1|0)&Co2[931]);

        Sum2[933]<=1^0^Co2[932];
        Co2[933]<=(1&0|(1|0)&Co2[932]);

        Sum2[934]<=1^0^Co2[933];
        Co2[934]<=(1&0|(1|0)&Co2[933]);

        Sum2[935]<=1^0^Co2[934];
        Co2[935]<=(1&0|(1|0)&Co2[934]);

        Sum2[936]<=1^0^Co2[935];
        Co2[936]<=(1&0|(1|0)&Co2[935]);

        Sum2[937]<=1^0^Co2[936];
        Co2[937]<=(1&0|(1|0)&Co2[936]);

        Sum2[938]<=1^0^Co2[937];
        Co2[938]<=(1&0|(1|0)&Co2[937]);

        Sum2[939]<=1^0^Co2[938];
        Co2[939]<=(1&0|(1|0)&Co2[938]);

        Sum2[940]<=1^0^Co2[939];
        Co2[940]<=(1&0|(1|0)&Co2[939]);

        Sum2[941]<=1^0^Co2[940];
        Co2[941]<=(1&0|(1|0)&Co2[940]);

        Sum2[942]<=1^0^Co2[941];
        Co2[942]<=(1&0|(1|0)&Co2[941]);

        Sum2[943]<=1^0^Co2[942];
        Co2[943]<=(1&0|(1|0)&Co2[942]);

        Sum2[944]<=1^0^Co2[943];
        Co2[944]<=(1&0|(1|0)&Co2[943]);

        Sum2[945]<=1^0^Co2[944];
        Co2[945]<=(1&0|(1|0)&Co2[944]);

        Sum2[946]<=1^0^Co2[945];
        Co2[946]<=(1&0|(1|0)&Co2[945]);

        Sum2[947]<=1^0^Co2[946];
        Co2[947]<=(1&0|(1|0)&Co2[946]);

        Sum2[948]<=1^0^Co2[947];
        Co2[948]<=(1&0|(1|0)&Co2[947]);

        Sum2[949]<=1^0^Co2[948];
        Co2[949]<=(1&0|(1|0)&Co2[948]);

        Sum2[950]<=1^0^Co2[949];
        Co2[950]<=(1&0|(1|0)&Co2[949]);

        Sum2[951]<=1^0^Co2[950];
        Co2[951]<=(1&0|(1|0)&Co2[950]);

        Sum2[952]<=1^0^Co2[951];
        Co2[952]<=(1&0|(1|0)&Co2[951]);

        Sum2[953]<=1^0^Co2[952];
        Co2[953]<=(1&0|(1|0)&Co2[952]);

        Sum2[954]<=1^0^Co2[953];
        Co2[954]<=(1&0|(1|0)&Co2[953]);

        Sum2[955]<=1^0^Co2[954];
        Co2[955]<=(1&0|(1|0)&Co2[954]);

        Sum2[956]<=1^0^Co2[955];
        Co2[956]<=(1&0|(1|0)&Co2[955]);

        Sum2[957]<=1^0^Co2[956];
        Co2[957]<=(1&0|(1|0)&Co2[956]);

        Sum2[958]<=1^0^Co2[957];
        Co2[958]<=(1&0|(1|0)&Co2[957]);

        Sum2[959]<=1^0^Co2[958];
        Co2[959]<=(1&0|(1|0)&Co2[958]);

        Sum2[960]<=1^0^Co2[959];
        Co2[960]<=(1&0|(1|0)&Co2[959]);

        Sum2[961]<=1^0^Co2[960];
        Co2[961]<=(1&0|(1|0)&Co2[960]);

        Sum2[962]<=1^0^Co2[961];
        Co2[962]<=(1&0|(1|0)&Co2[961]);

        Sum2[963]<=1^0^Co2[962];
        Co2[963]<=(1&0|(1|0)&Co2[962]);

        Sum2[964]<=1^0^Co2[963];
        Co2[964]<=(1&0|(1|0)&Co2[963]);

        Sum2[965]<=1^0^Co2[964];
        Co2[965]<=(1&0|(1|0)&Co2[964]);

        Sum2[966]<=1^0^Co2[965];
        Co2[966]<=(1&0|(1|0)&Co2[965]);

        Sum2[967]<=1^0^Co2[966];
        Co2[967]<=(1&0|(1|0)&Co2[966]);

        Sum2[968]<=1^0^Co2[967];
        Co2[968]<=(1&0|(1|0)&Co2[967]);

        Sum2[969]<=1^0^Co2[968];
        Co2[969]<=(1&0|(1|0)&Co2[968]);

        Sum2[970]<=1^0^Co2[969];
        Co2[970]<=(1&0|(1|0)&Co2[969]);

        Sum2[971]<=1^0^Co2[970];
        Co2[971]<=(1&0|(1|0)&Co2[970]);

        Sum2[972]<=1^0^Co2[971];
        Co2[972]<=(1&0|(1|0)&Co2[971]);

        Sum2[973]<=1^0^Co2[972];
        Co2[973]<=(1&0|(1|0)&Co2[972]);

        Sum2[974]<=1^0^Co2[973];
        Co2[974]<=(1&0|(1|0)&Co2[973]);

        Sum2[975]<=1^0^Co2[974];
        Co2[975]<=(1&0|(1|0)&Co2[974]);

        Sum2[976]<=1^0^Co2[975];
        Co2[976]<=(1&0|(1|0)&Co2[975]);

        Sum2[977]<=1^0^Co2[976];
        Co2[977]<=(1&0|(1|0)&Co2[976]);

        Sum2[978]<=1^0^Co2[977];
        Co2[978]<=(1&0|(1|0)&Co2[977]);

        Sum2[979]<=1^0^Co2[978];
        Co2[979]<=(1&0|(1|0)&Co2[978]);

        Sum2[980]<=1^0^Co2[979];
        Co2[980]<=(1&0|(1|0)&Co2[979]);

        Sum2[981]<=1^0^Co2[980];
        Co2[981]<=(1&0|(1|0)&Co2[980]);

        Sum2[982]<=1^0^Co2[981];
        Co2[982]<=(1&0|(1|0)&Co2[981]);

        Sum2[983]<=1^0^Co2[982];
        Co2[983]<=(1&0|(1|0)&Co2[982]);

        Sum2[984]<=1^0^Co2[983];
        Co2[984]<=(1&0|(1|0)&Co2[983]);

        Sum2[985]<=1^0^Co2[984];
        Co2[985]<=(1&0|(1|0)&Co2[984]);

        Sum2[986]<=1^0^Co2[985];
        Co2[986]<=(1&0|(1|0)&Co2[985]);

        Sum2[987]<=1^0^Co2[986];
        Co2[987]<=(1&0|(1|0)&Co2[986]);

        Sum2[988]<=1^0^Co2[987];
        Co2[988]<=(1&0|(1|0)&Co2[987]);

        Sum2[989]<=1^0^Co2[988];
        Co2[989]<=(1&0|(1|0)&Co2[988]);

        Sum2[990]<=1^0^Co2[989];
        Co2[990]<=(1&0|(1|0)&Co2[989]);

        Sum2[991]<=1^0^Co2[990];
        Co2[991]<=(1&0|(1|0)&Co2[990]);

        Sum2[992]<=1^0^Co2[991];
        Co2[992]<=(1&0|(1|0)&Co2[991]);

        Sum2[993]<=1^0^Co2[992];
        Co2[993]<=(1&0|(1|0)&Co2[992]);

        Sum2[994]<=1^0^Co2[993];
        Co2[994]<=(1&0|(1|0)&Co2[993]);

        Sum2[995]<=1^0^Co2[994];
        Co2[995]<=(1&0|(1|0)&Co2[994]);

        Sum2[996]<=1^0^Co2[995];
        Co2[996]<=(1&0|(1|0)&Co2[995]);

        Sum2[997]<=1^0^Co2[996];
        Co2[997]<=(1&0|(1|0)&Co2[996]);

        Sum2[998]<=1^0^Co2[997];
        Co2[998]<=(1&0|(1|0)&Co2[997]);

        Sum2[999]<=1^0^Co2[998];
        Co2[999]<=(1&0|(1|0)&Co2[998]);

        Sum2[1000]<=1^0^Co2[999];
        Co2[1000]<=(1&0|(1|0)&Co2[999]);

        Sum2[1001]<=1^0^Co2[1000];
        Co2[1001]<=(1&0|(1|0)&Co2[1000]);

        Sum2[1002]<=1^0^Co2[1001];
        Co2[1002]<=(1&0|(1|0)&Co2[1001]);

        Sum2[1003]<=1^0^Co2[1002];
        Co2[1003]<=(1&0|(1|0)&Co2[1002]);

        Sum2[1004]<=1^0^Co2[1003];
        Co2[1004]<=(1&0|(1|0)&Co2[1003]);

        Sum2[1005]<=1^0^Co2[1004];
        Co2[1005]<=(1&0|(1|0)&Co2[1004]);

        Sum2[1006]<=1^0^Co2[1005];
        Co2[1006]<=(1&0|(1|0)&Co2[1005]);

        Sum2[1007]<=1^0^Co2[1006];
        Co2[1007]<=(1&0|(1|0)&Co2[1006]);

        Sum2[1008]<=1^0^Co2[1007];
        Co2[1008]<=(1&0|(1|0)&Co2[1007]);

        Sum2[1009]<=1^0^Co2[1008];
        Co2[1009]<=(1&0|(1|0)&Co2[1008]);

        Sum2[1010]<=1^0^Co2[1009];
        Co2[1010]<=(1&0|(1|0)&Co2[1009]);

        Sum2[1011]<=1^0^Co2[1010];
        Co2[1011]<=(1&0|(1|0)&Co2[1010]);

        Sum2[1012]<=1^0^Co2[1011];
        Co2[1012]<=(1&0|(1|0)&Co2[1011]);

        Sum2[1013]<=1^0^Co2[1012];
        Co2[1013]<=(1&0|(1|0)&Co2[1012]);

        Sum2[1014]<=1^0^Co2[1013];
        Co2[1014]<=(1&0|(1|0)&Co2[1013]);

        Sum2[1015]<=1^0^Co2[1014];
        Co2[1015]<=(1&0|(1|0)&Co2[1014]);

        Sum2[1016]<=1^0^Co2[1015];
        Co2[1016]<=(1&0|(1|0)&Co2[1015]);

        Sum2[1017]<=1^0^Co2[1016];
        Co2[1017]<=(1&0|(1|0)&Co2[1016]);

        Sum2[1018]<=1^0^Co2[1017];
        Co2[1018]<=(1&0|(1|0)&Co2[1017]);

        Sum2[1019]<=1^0^Co2[1018];
        Co2[1019]<=(1&0|(1|0)&Co2[1018]);

        Sum2[1020]<=1^0^Co2[1019];
        Co2[1020]<=(1&0|(1|0)&Co2[1019]);

        Sum2[1021]<=1^0^Co2[1020];
        Co2[1021]<=(1&0|(1|0)&Co2[1020]);

        Sum2[1022]<=1^0^Co2[1021];
        Co2[1022]<=(1&0|(1|0)&Co2[1021]);

        Sum2[1023]<=1^0^Co2[1022];
        Co2[1023]<=(1&0|(1|0)&Co2[1022]);
        */
end

//assign out_data = Sum2;
assign Out = Co2[1023];

endmodule
